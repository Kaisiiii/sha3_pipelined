module pad (
    input [1087:0] data_in,
    input [10:0] data_length,
    output reg [1087:0] data_out,
    output reg [1087:0] data_next
);

    always@(*) begin
        if ((data_length >= 0) && (data_length <= 1088)) begin
				//data_out = 'd0;
            if (data_length == 0) begin
                data_out = 1088'h1f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
                data_next = 1088'b0;
            end else if (data_length == 1088) begin
                data_out = data_in;
                data_next = 1088'h1f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else if (data_length == 1087) begin
                data_out = {data_in[1087:8], 1'h1, data_in[7:1]};
                data_next = 1088'h0f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else if (data_length == 1086) begin
                data_out = {data_in[1087:8], 2'h3, data_in[7:2]};
                data_next = 1088'h07000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else if (data_length == 1085) begin
                data_out = {data_in[1087:8], 3'h7, data_in[7:3]};
                data_next = 1088'h03000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else if (data_length == 1084) begin
                data_out = {data_in[1087:8], 4'hf, data_in[7:4]};
                data_next = 1088'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else if (data_length == 1083) begin
                data_out = {data_in[1087:8], 5'h1f, data_in[7:5]};
                data_next = 1088'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080;
            end else begin
                case (data_length)
                    1   : data_out = {                    7'h1f, data_in[1087],             {1072{1'b0}}, 8'h80};
                    2   : data_out = {                    6'h1f, data_in[1087:1086],        {1072{1'b0}}, 8'h80};
                    3   : data_out = {                    5'h1f, data_in[1087:1085],        {1072{1'b0}}, 8'h80};
                    4   : data_out = {                    4'hf,  data_in[1087:1084], 8'h1,  {1064{1'b0}}, 8'h80};
                    5   : data_out = {                    3'h7,  data_in[1087:1083], 8'h3,  {1064{1'b0}}, 8'h80};
                    6   : data_out = {                    2'h3,  data_in[1087:1082], 8'h7,  {1064{1'b0}}, 8'h80};
                    7   : data_out = {                    1'h1,  data_in[1087:1081], 8'hf,  {1064{1'b0}}, 8'h80};
                    8   : data_out = {data_in[1087:1080],                            8'h1f, {1064{1'b0}}, 8'h80};
                    
                    9   : data_out = {data_in[1087:1080], 7'h1f, data_in[1079],             {1064{1'b0}}, 8'h80};
                    10  : data_out = {data_in[1087:1080], 6'h1f, data_in[1079:1078],        {1064{1'b0}}, 8'h80};
                    11  : data_out = {data_in[1087:1080], 5'h1f, data_in[1079:1077],        {1064{1'b0}}, 8'h80};
                    12  : data_out = {data_in[1087:1080], 4'hf,  data_in[1079:1076], 8'h1,  {1056{1'b0}}, 8'h80};
                    13  : data_out = {data_in[1087:1080], 3'h7,  data_in[1079:1075], 8'h3,  {1056{1'b0}}, 8'h80};
                    14  : data_out = {data_in[1087:1080], 2'h3,  data_in[1079:1074], 8'h7,  {1056{1'b0}}, 8'h80};
                    15  : data_out = {data_in[1087:1080], 1'h1,  data_in[1079:1073], 8'hf,  {1056{1'b0}}, 8'h80};
                    16  : data_out = {data_in[1087:1072],                            8'h1f, {1056{1'b0}}, 8'h80};
                    
                    17  : data_out = {data_in[1087:1072], 7'h1f, data_in[1071],             {1056{1'b0}}, 8'h80};
                    18  : data_out = {data_in[1087:1072], 6'h1f, data_in[1071:1070],        {1056{1'b0}}, 8'h80};
                    19  : data_out = {data_in[1087:1072], 5'h1f, data_in[1071:1069],        {1056{1'b0}}, 8'h80};
                    20  : data_out = {data_in[1087:1072], 4'hf,  data_in[1071:1068], 8'h1,  {1048{1'b0}}, 8'h80};
                    21  : data_out = {data_in[1087:1072], 3'h7,  data_in[1071:1067], 8'h3,  {1048{1'b0}}, 8'h80};
                    22  : data_out = {data_in[1087:1072], 2'h3,  data_in[1071:1066], 8'h7,  {1048{1'b0}}, 8'h80};
                    23  : data_out = {data_in[1087:1072], 1'h1,  data_in[1071:1065], 8'hf,  {1048{1'b0}}, 8'h80};
                    24  : data_out = {data_in[1087:1064],                            8'h1f, {1048{1'b0}}, 8'h80};
                    
                    25  : data_out = {data_in[1087:1064], 7'h1f, data_in[1063],             {1048{1'b0}}, 8'h80};
                    26  : data_out = {data_in[1087:1064], 6'h1f, data_in[1063:1062],        {1048{1'b0}}, 8'h80};
                    27  : data_out = {data_in[1087:1064], 5'h1f, data_in[1063:1061],        {1048{1'b0}}, 8'h80};
                    28  : data_out = {data_in[1087:1064], 4'hf,  data_in[1063:1060], 8'h1,  {1040{1'b0}}, 8'h80};
                    29  : data_out = {data_in[1087:1064], 3'h7,  data_in[1063:1059], 8'h3,  {1040{1'b0}}, 8'h80};
                    30  : data_out = {data_in[1087:1064], 2'h3,  data_in[1063:1058], 8'h7,  {1040{1'b0}}, 8'h80};
                    31  : data_out = {data_in[1087:1064], 1'h1,  data_in[1063:1057], 8'hf,  {1040{1'b0}}, 8'h80};
                    32  : data_out = {data_in[1087:1056],                            8'h1f, {1040{1'b0}}, 8'h80};
                    
                    33  : data_out = {data_in[1087:1056], 7'h1f, data_in[1055],             {1040{1'b0}}, 8'h80};
                    34  : data_out = {data_in[1087:1056], 6'h1f, data_in[1055:1054],        {1040{1'b0}}, 8'h80};
                    35  : data_out = {data_in[1087:1056], 5'h1f, data_in[1055:1053],        {1040{1'b0}}, 8'h80};
                    36  : data_out = {data_in[1087:1056], 4'hf,  data_in[1055:1052], 8'h1,  {1032{1'b0}}, 8'h80};
                    37  : data_out = {data_in[1087:1056], 3'h7,  data_in[1055:1051], 8'h3,  {1032{1'b0}}, 8'h80};
                    38  : data_out = {data_in[1087:1056], 2'h3,  data_in[1055:1050], 8'h7,  {1032{1'b0}}, 8'h80};
                    39  : data_out = {data_in[1087:1056], 1'h1,  data_in[1055:1049], 8'hf,  {1032{1'b0}}, 8'h80};
                    40  : data_out = {data_in[1087:1048],                            8'h1f, {1032{1'b0}}, 8'h80};
                    
                    41  : data_out = {data_in[1087:1048], 7'h1f, data_in[1047],             {1032{1'b0}}, 8'h80};
                    42  : data_out = {data_in[1087:1048], 6'h1f, data_in[1047:1046],        {1032{1'b0}}, 8'h80};
                    43  : data_out = {data_in[1087:1048], 5'h1f, data_in[1047:1045],        {1032{1'b0}}, 8'h80};
                    44  : data_out = {data_in[1087:1048], 4'hf,  data_in[1047:1044], 8'h1,  {1024{1'b0}}, 8'h80};
                    45  : data_out = {data_in[1087:1048], 3'h7,  data_in[1047:1043], 8'h3,  {1024{1'b0}}, 8'h80};
                    46  : data_out = {data_in[1087:1048], 2'h3,  data_in[1047:1042], 8'h7,  {1024{1'b0}}, 8'h80};
                    47  : data_out = {data_in[1087:1048], 1'h1,  data_in[1047:1041], 8'hf,  {1024{1'b0}}, 8'h80};
                    48  : data_out = {data_in[1087:1040],                            8'h1f, {1024{1'b0}}, 8'h80};
                    
                    49  : data_out = {data_in[1087:1040], 7'h1f, data_in[1039],             {1024{1'b0}}, 8'h80};
                    50  : data_out = {data_in[1087:1040], 6'h1f, data_in[1039:1038],        {1024{1'b0}}, 8'h80};
                    51  : data_out = {data_in[1087:1040], 5'h1f, data_in[1039:1037],        {1024{1'b0}}, 8'h80};
                    52  : data_out = {data_in[1087:1040], 4'hf,  data_in[1039:1036], 8'h1,  {1016{1'b0}}, 8'h80};
                    53  : data_out = {data_in[1087:1040], 3'h7,  data_in[1039:1035], 8'h3,  {1016{1'b0}}, 8'h80};
                    54  : data_out = {data_in[1087:1040], 2'h3,  data_in[1039:1034], 8'h7,  {1016{1'b0}}, 8'h80};
                    55  : data_out = {data_in[1087:1040], 1'h1,  data_in[1039:1033], 8'hf,  {1016{1'b0}}, 8'h80};
                    56  : data_out = {data_in[1087:1032],                            8'h1f, {1016{1'b0}}, 8'h80};
                    
                    57  : data_out = {data_in[1087:1032], 7'h1f, data_in[1031],             {1016{1'b0}}, 8'h80};
                    58  : data_out = {data_in[1087:1032], 6'h1f, data_in[1031:1030],        {1016{1'b0}}, 8'h80};
                    59  : data_out = {data_in[1087:1032], 5'h1f, data_in[1031:1029],        {1016{1'b0}}, 8'h80};
                    60  : data_out = {data_in[1087:1032], 4'hf,  data_in[1031:1028], 8'h1,  {1008{1'b0}}, 8'h80};
                    61  : data_out = {data_in[1087:1032], 3'h7,  data_in[1031:1027], 8'h3,  {1008{1'b0}}, 8'h80};
                    62  : data_out = {data_in[1087:1032], 2'h3,  data_in[1031:1026], 8'h7,  {1008{1'b0}}, 8'h80};
                    63  : data_out = {data_in[1087:1032], 1'h1,  data_in[1031:1025], 8'hf,  {1008{1'b0}}, 8'h80};
                    64  : data_out = {data_in[1087:1024],                            8'h1f, {1008{1'b0}}, 8'h80};
                    
                    65  : data_out = {data_in[1087:1024], 7'h1f, data_in[1023],             {1008{1'b0}}, 8'h80};
                    66  : data_out = {data_in[1087:1024], 6'h1f, data_in[1023:1022],        {1008{1'b0}}, 8'h80};
                    67  : data_out = {data_in[1087:1024], 5'h1f, data_in[1023:1021],        {1008{1'b0}}, 8'h80};
                    68  : data_out = {data_in[1087:1024], 4'hf,  data_in[1023:1020], 8'h1,  {1000{1'b0}}, 8'h80};
                    69  : data_out = {data_in[1087:1024], 3'h7,  data_in[1023:1019], 8'h3,  {1000{1'b0}}, 8'h80};
                    70  : data_out = {data_in[1087:1024], 2'h3,  data_in[1023:1018], 8'h7,  {1000{1'b0}}, 8'h80};
                    71  : data_out = {data_in[1087:1024], 1'h1,  data_in[1023:1017], 8'hf,  {1000{1'b0}}, 8'h80};
                    72  : data_out = {data_in[1087:1016],                            8'h1f, {1000{1'b0}}, 8'h80};
                    
                    73  : data_out = {data_in[1087:1016], 7'h1f, data_in[1015],             {1000{1'b0}}, 8'h80};
                    74  : data_out = {data_in[1087:1016], 6'h1f, data_in[1015:1014],        {1000{1'b0}}, 8'h80};
                    75  : data_out = {data_in[1087:1016], 5'h1f, data_in[1015:1013],        {1000{1'b0}}, 8'h80};
                    76  : data_out = {data_in[1087:1016], 4'hf,  data_in[1015:1012], 8'h1,  {992{1'b0}},  8'h80};
                    77  : data_out = {data_in[1087:1016], 3'h7,  data_in[1015:1011], 8'h3,  {992{1'b0}},  8'h80};
                    78  : data_out = {data_in[1087:1016], 2'h3,  data_in[1015:1010], 8'h7,  {992{1'b0}},  8'h80};
                    79  : data_out = {data_in[1087:1016], 1'h1,  data_in[1015:1009], 8'hf,  {992{1'b0}},  8'h80};
                    80  : data_out = {data_in[1087:1008],                            8'h1f, {992{1'b0}},  8'h80};
                    
                    81  : data_out = {data_in[1087:1008], 7'h1f, data_in[1007],             {992{1'b0}},  8'h80};
                    82  : data_out = {data_in[1087:1008], 6'h1f, data_in[1007:1006],        {992{1'b0}},  8'h80};
                    83  : data_out = {data_in[1087:1008], 5'h1f, data_in[1007:1005],        {992{1'b0}},  8'h80};
                    84  : data_out = {data_in[1087:1008], 4'hf,  data_in[1007:1004], 8'h1,  {984{1'b0}},  8'h80};
                    85  : data_out = {data_in[1087:1008], 3'h7,  data_in[1007:1003], 8'h3,  {984{1'b0}},  8'h80};
                    86  : data_out = {data_in[1087:1008], 2'h3,  data_in[1007:1002], 8'h7,  {984{1'b0}},  8'h80};
                    87  : data_out = {data_in[1087:1008], 1'h1,  data_in[1007:1001], 8'hf,  {984{1'b0}},  8'h80};
                    88  : data_out = {data_in[1087:1000],                            8'h1f, {984{1'b0}},  8'h80};
                    
                    89  : data_out = {data_in[1087:1000], 7'h1f, data_in[999],              {984{1'b0}},  8'h80};
                    90  : data_out = {data_in[1087:1000], 6'h1f, data_in[999:998],          {984{1'b0}},  8'h80};
                    91  : data_out = {data_in[1087:1000], 5'h1f, data_in[999:997],          {984{1'b0}},  8'h80};
                    92  : data_out = {data_in[1087:1000], 4'hf,  data_in[999:996],   8'h1,  {976{1'b0}},  8'h80};
                    93  : data_out = {data_in[1087:1000], 3'h7,  data_in[999:995],   8'h3,  {976{1'b0}},  8'h80};
                    94  : data_out = {data_in[1087:1000], 2'h3,  data_in[999:994],   8'h7,  {976{1'b0}},  8'h80};
                    95  : data_out = {data_in[1087:1000], 1'h1,  data_in[999:993],   8'hf,  {976{1'b0}},  8'h80};
                    96  : data_out = {data_in[1087:992],                             8'h1f, {976{1'b0}},  8'h80};
                    
                    97  : data_out = {data_in[1087:992],  7'h1f, data_in[991],              {976{1'b0}},  8'h80};
                    98  : data_out = {data_in[1087:992],  6'h1f, data_in[991:990],          {976{1'b0}},  8'h80};
                    99  : data_out = {data_in[1087:992],  5'h1f, data_in[991:989],          {976{1'b0}},  8'h80};
                    100 : data_out = {data_in[1087:992],  4'hf,  data_in[991:988],   8'h1,  {968{1'b0}},  8'h80};
                    101 : data_out = {data_in[1087:992],  3'h7,  data_in[991:987],   8'h3,  {968{1'b0}},  8'h80};
                    102 : data_out = {data_in[1087:992],  2'h3,  data_in[991:986],   8'h7,  {968{1'b0}},  8'h80};
                    103 : data_out = {data_in[1087:992],  1'h1,  data_in[991:985],   8'hf,  {968{1'b0}},  8'h80};
                    104 : data_out = {data_in[1087:984],                             8'h1f, {968{1'b0}},  8'h80};
                    
                    105 : data_out = {data_in[1087:984],  7'h1f, data_in[983],              {968{1'b0}},  8'h80};
                    106 : data_out = {data_in[1087:984],  6'h1f, data_in[983:982],          {968{1'b0}},  8'h80};
                    107 : data_out = {data_in[1087:984],  5'h1f, data_in[983:981],          {968{1'b0}},  8'h80};
                    108 : data_out = {data_in[1087:984],  4'hf,  data_in[983:980],   8'h1,  {960{1'b0}},  8'h80};
                    109 : data_out = {data_in[1087:984],  3'h7,  data_in[983:979],   8'h3,  {960{1'b0}},  8'h80};
                    110 : data_out = {data_in[1087:984],  2'h3,  data_in[983:978],   8'h7,  {960{1'b0}},  8'h80};
                    111 : data_out = {data_in[1087:984],  1'h1,  data_in[983:977],   8'hf,  {960{1'b0}},  8'h80};
                    112 : data_out = {data_in[1087:976],                             8'h1f, {960{1'b0}},  8'h80};

                    113 : data_out = {data_in[1087:976],  7'h1f, data_in[975],              {960{1'b0}},  8'h80};
                    114 : data_out = {data_in[1087:976],  6'h1f, data_in[975:974],          {960{1'b0}},  8'h80};
                    115 : data_out = {data_in[1087:976],  5'h1f, data_in[975:973],          {960{1'b0}},  8'h80};
                    116 : data_out = {data_in[1087:976],  4'hf,  data_in[975:972],   8'h1,  {952{1'b0}},  8'h80};
                    117 : data_out = {data_in[1087:976],  3'h7,  data_in[975:971],   8'h3,  {952{1'b0}},  8'h80};
                    118 : data_out = {data_in[1087:976],  2'h3,  data_in[975:970],   8'h7,  {952{1'b0}},  8'h80};
                    119 : data_out = {data_in[1087:976],  1'h1,  data_in[975:969],   8'hf,  {952{1'b0}},  8'h80};
                    120 : data_out = {data_in[1087:968],                             8'h1f, {952{1'b0}},  8'h80};

                    121 : data_out = {data_in[1087:968],  7'h1f, data_in[967],              {952{1'b0}},  8'h80};
                    122 : data_out = {data_in[1087:968],  6'h1f, data_in[967:966],          {952{1'b0}},  8'h80};
                    123 : data_out = {data_in[1087:968],  5'h1f, data_in[967:965],          {952{1'b0}},  8'h80};
                    124 : data_out = {data_in[1087:968],  4'hf,  data_in[967:964],   8'h1,  {944{1'b0}},  8'h80};
                    125 : data_out = {data_in[1087:968],  3'h7,  data_in[967:963],   8'h3,  {944{1'b0}},  8'h80};
                    126 : data_out = {data_in[1087:968],  2'h3,  data_in[967:962],   8'h7,  {944{1'b0}},  8'h80};
                    127 : data_out = {data_in[1087:968],  1'h1,  data_in[967:961],   8'hf,  {944{1'b0}},  8'h80};
                    128 : data_out = {data_in[1087:960],                             8'h1f, {944{1'b0}},  8'h80};

                    129 : data_out = {data_in[1087:960],  7'h1f, data_in[959],              {944{1'b0}},  8'h80};
                    130 : data_out = {data_in[1087:960],  6'h1f, data_in[959:958],          {944{1'b0}},  8'h80};
                    131 : data_out = {data_in[1087:960],  5'h1f, data_in[959:957],          {944{1'b0}},  8'h80};
                    132 : data_out = {data_in[1087:960],  4'hf,  data_in[959:956],   8'h1,  {936{1'b0}},  8'h80};
                    133 : data_out = {data_in[1087:960],  3'h7,  data_in[959:955],   8'h3,  {936{1'b0}},  8'h80};
                    134 : data_out = {data_in[1087:960],  2'h3,  data_in[959:954],   8'h7,  {936{1'b0}},  8'h80};
                    135 : data_out = {data_in[1087:960],  1'h1,  data_in[959:953],   8'hf,  {936{1'b0}},  8'h80};
                    136 : data_out = {data_in[1087:952],                             8'h1f, {936{1'b0}},  8'h80};

                    137 : data_out = {data_in[1087:952],  7'h1f, data_in[951],              {936{1'b0}},  8'h80};
                    138 : data_out = {data_in[1087:952],  6'h1f, data_in[951:950],          {936{1'b0}},  8'h80};
                    139 : data_out = {data_in[1087:952],  5'h1f, data_in[951:949],          {936{1'b0}},  8'h80};
                    140 : data_out = {data_in[1087:952],  4'hf,  data_in[951:948],   8'h1,  {928{1'b0}},  8'h80};
                    141 : data_out = {data_in[1087:952],  3'h7,  data_in[951:947],   8'h3,  {928{1'b0}},  8'h80};
                    142 : data_out = {data_in[1087:952],  2'h3,  data_in[951:946],   8'h7,  {928{1'b0}},  8'h80};
                    143 : data_out = {data_in[1087:952],  1'h1,  data_in[951:945],   8'hf,  {928{1'b0}},  8'h80};
                    144 : data_out = {data_in[1087:944],                             8'h1f, {928{1'b0}},  8'h80};

                    145 : data_out = {data_in[1087:944],  7'h1f, data_in[943],              {928{1'b0}},  8'h80};
                    146 : data_out = {data_in[1087:944],  6'h1f, data_in[943:942],          {928{1'b0}},  8'h80};
                    147 : data_out = {data_in[1087:944],  5'h1f, data_in[943:941],          {928{1'b0}},  8'h80};
                    148 : data_out = {data_in[1087:944],  4'hf,  data_in[943:940],   8'h1,  {920{1'b0}},  8'h80};
                    149 : data_out = {data_in[1087:944],  3'h7,  data_in[943:939],   8'h3,  {920{1'b0}},  8'h80};
                    150 : data_out = {data_in[1087:944],  2'h3,  data_in[943:938],   8'h7,  {920{1'b0}},  8'h80};
                    151 : data_out = {data_in[1087:944],  1'h1,  data_in[943:937],   8'hf,  {920{1'b0}},  8'h80};
                    152 : data_out = {data_in[1087:936],                             8'h1f, {920{1'b0}},  8'h80};

                    153 : data_out = {data_in[1087:936],  7'h1f, data_in[935],              {920{1'b0}},  8'h80};
                    154 : data_out = {data_in[1087:936],  6'h1f, data_in[935:934],          {920{1'b0}},  8'h80};
                    155 : data_out = {data_in[1087:936],  5'h1f, data_in[935:933],          {920{1'b0}},  8'h80};
                    156 : data_out = {data_in[1087:936],  4'hf,  data_in[935:932],   8'h1,  {912{1'b0}},  8'h80};
                    157 : data_out = {data_in[1087:936],  3'h7,  data_in[935:931],   8'h3,  {912{1'b0}},  8'h80};
                    158 : data_out = {data_in[1087:936],  2'h3,  data_in[935:930],   8'h7,  {912{1'b0}},  8'h80};
                    159 : data_out = {data_in[1087:936],  1'h1,  data_in[935:929],   8'hf,  {912{1'b0}},  8'h80};
                    160 : data_out = {data_in[1087:928],                             8'h1f, {912{1'b0}},  8'h80};

                    161 : data_out = {data_in[1087:928],  7'h1f, data_in[927],              {912{1'b0}},  8'h80};
                    162 : data_out = {data_in[1087:928],  6'h1f, data_in[927:926],          {912{1'b0}},  8'h80};
                    163 : data_out = {data_in[1087:928],  5'h1f, data_in[927:925],          {912{1'b0}},  8'h80};
                    164 : data_out = {data_in[1087:928],  4'hf,  data_in[927:924],   8'h1,  {904{1'b0}},  8'h80};
                    165 : data_out = {data_in[1087:928],  3'h7,  data_in[927:923],   8'h3,  {904{1'b0}},  8'h80};
                    166 : data_out = {data_in[1087:928],  2'h3,  data_in[927:922],   8'h7,  {904{1'b0}},  8'h80};
                    167 : data_out = {data_in[1087:928],  1'h1,  data_in[927:921],   8'hf,  {904{1'b0}},  8'h80};
                    168 : data_out = {data_in[1087:920],                             8'h1f, {904{1'b0}},  8'h80};

                    169 : data_out = {data_in[1087:920],  7'h1f, data_in[919],              {904{1'b0}},  8'h80};
                    170 : data_out = {data_in[1087:920],  6'h1f, data_in[919:918],          {904{1'b0}},  8'h80};
                    171 : data_out = {data_in[1087:920],  5'h1f, data_in[919:917],          {904{1'b0}},  8'h80};
                    172 : data_out = {data_in[1087:920],  4'hf,  data_in[919:916],   8'h1,  {896{1'b0}},  8'h80};
                    173 : data_out = {data_in[1087:920],  3'h7,  data_in[919:915],   8'h3,  {896{1'b0}},  8'h80};
                    174 : data_out = {data_in[1087:920],  2'h3,  data_in[919:914],   8'h7,  {896{1'b0}},  8'h80};
                    175 : data_out = {data_in[1087:920],  1'h1,  data_in[919:913],   8'hf,  {896{1'b0}},  8'h80};
                    176 : data_out = {data_in[1087:912],                             8'h1f, {896{1'b0}},  8'h80};

                    177 : data_out = {data_in[1087:912],  7'h1f, data_in[911],              {896{1'b0}},  8'h80};
                    178 : data_out = {data_in[1087:912],  6'h1f, data_in[911:910],          {896{1'b0}},  8'h80};
                    179 : data_out = {data_in[1087:912],  5'h1f, data_in[911:909],          {896{1'b0}},  8'h80};
                    180 : data_out = {data_in[1087:912],  4'hf,  data_in[911:908],   8'h1,  {888{1'b0}},  8'h80};
                    181 : data_out = {data_in[1087:912],  3'h7,  data_in[911:907],   8'h3,  {888{1'b0}},  8'h80};
                    182 : data_out = {data_in[1087:912],  2'h3,  data_in[911:906],   8'h7,  {888{1'b0}},  8'h80};
                    183 : data_out = {data_in[1087:912],  1'h1,  data_in[911:905],   8'hf,  {888{1'b0}},  8'h80};
                    184 : data_out = {data_in[1087:904],                             8'h1f, {888{1'b0}},  8'h80};

                    185 : data_out = {data_in[1087:904],  7'h1f, data_in[903],              {888{1'b0}},  8'h80};
                    186 : data_out = {data_in[1087:904],  6'h1f, data_in[903:902],          {888{1'b0}},  8'h80};
                    187 : data_out = {data_in[1087:904],  5'h1f, data_in[903:901],          {888{1'b0}},  8'h80};
                    188 : data_out = {data_in[1087:904],  4'hf,  data_in[903:900],   8'h1,  {880{1'b0}},  8'h80};
                    189 : data_out = {data_in[1087:904],  3'h7,  data_in[903:899],   8'h3,  {880{1'b0}},  8'h80};
                    190 : data_out = {data_in[1087:904],  2'h3,  data_in[903:898],   8'h7,  {880{1'b0}},  8'h80};
                    191 : data_out = {data_in[1087:904],  1'h1,  data_in[903:897],   8'hf,  {880{1'b0}},  8'h80};
                    192 : data_out = {data_in[1087:896],                             8'h1f, {880{1'b0}},  8'h80};

                    193 : data_out = {data_in[1087:896],  7'h1f, data_in[895],              {880{1'b0}},  8'h80};
                    194 : data_out = {data_in[1087:896],  6'h1f, data_in[895:894],          {880{1'b0}},  8'h80};
                    195 : data_out = {data_in[1087:896],  5'h1f, data_in[895:893],          {880{1'b0}},  8'h80};
                    196 : data_out = {data_in[1087:896],  4'hf,  data_in[895:892],   8'h1,  {872{1'b0}},  8'h80};
                    197 : data_out = {data_in[1087:896],  3'h7,  data_in[895:891],   8'h3,  {872{1'b0}},  8'h80};
                    198 : data_out = {data_in[1087:896],  2'h3,  data_in[895:890],   8'h7,  {872{1'b0}},  8'h80};
                    199 : data_out = {data_in[1087:896],  1'h1,  data_in[895:889],   8'hf,  {872{1'b0}},  8'h80};
                    200 : data_out = {data_in[1087:888],                             8'h1f, {872{1'b0}},  8'h80};

                    201 : data_out = {data_in[1087:888],  7'h1f, data_in[887],              {872{1'b0}},  8'h80};
                    202 : data_out = {data_in[1087:888],  6'h1f, data_in[887:886],          {872{1'b0}},  8'h80};
                    203 : data_out = {data_in[1087:888],  5'h1f, data_in[887:885],          {872{1'b0}},  8'h80};
                    204 : data_out = {data_in[1087:888],  4'hf,  data_in[887:884],   8'h1,  {864{1'b0}},  8'h80};
                    205 : data_out = {data_in[1087:888],  3'h7,  data_in[887:883],   8'h3,  {864{1'b0}},  8'h80};
                    206 : data_out = {data_in[1087:888],  2'h3,  data_in[887:882],   8'h7,  {864{1'b0}},  8'h80};
                    207 : data_out = {data_in[1087:888],  1'h1,  data_in[887:881],   8'hf,  {864{1'b0}},  8'h80};
                    208 : data_out = {data_in[1087:880],                             8'h1f, {864{1'b0}},  8'h80};

                    209 : data_out = {data_in[1087:880],  7'h1f, data_in[879],              {864{1'b0}},  8'h80};
                    210 : data_out = {data_in[1087:880],  6'h1f, data_in[879:878],          {864{1'b0}},  8'h80};
                    211 : data_out = {data_in[1087:880],  5'h1f, data_in[879:877],          {864{1'b0}},  8'h80};
                    212 : data_out = {data_in[1087:880],  4'hf,  data_in[879:876],   8'h1,  {856{1'b0}},  8'h80};
                    213 : data_out = {data_in[1087:880],  3'h7,  data_in[879:875],   8'h3,  {856{1'b0}},  8'h80};
                    214 : data_out = {data_in[1087:880],  2'h3,  data_in[879:874],   8'h7,  {856{1'b0}},  8'h80};
                    215 : data_out = {data_in[1087:880],  1'h1,  data_in[879:873],   8'hf,  {856{1'b0}},  8'h80};
                    216 : data_out = {data_in[1087:872],                             8'h1f, {856{1'b0}},  8'h80};

                    217 : data_out = {data_in[1087:872],  7'h1f, data_in[871],              {856{1'b0}},  8'h80};
                    218 : data_out = {data_in[1087:872],  6'h1f, data_in[871:870],          {856{1'b0}},  8'h80};
                    219 : data_out = {data_in[1087:872],  5'h1f, data_in[871:869],          {856{1'b0}},  8'h80};
                    220 : data_out = {data_in[1087:872],  4'hf,  data_in[871:868],   8'h1,  {848{1'b0}},  8'h80};
                    221 : data_out = {data_in[1087:872],  3'h7,  data_in[871:867],   8'h3,  {848{1'b0}},  8'h80};
                    222 : data_out = {data_in[1087:872],  2'h3,  data_in[871:866],   8'h7,  {848{1'b0}},  8'h80};
                    223 : data_out = {data_in[1087:872],  1'h1,  data_in[871:865],   8'hf,  {848{1'b0}},  8'h80};
                    224 : data_out = {data_in[1087:864],                             8'h1f, {848{1'b0}},  8'h80};

                    225 : data_out = {data_in[1087:864],  7'h1f, data_in[863],              {848{1'b0}},  8'h80};
                    226 : data_out = {data_in[1087:864],  6'h1f, data_in[863:862],          {848{1'b0}},  8'h80};
                    227 : data_out = {data_in[1087:864],  5'h1f, data_in[863:861],          {848{1'b0}},  8'h80};
                    228 : data_out = {data_in[1087:864],  4'hf,  data_in[863:860],   8'h1,  {840{1'b0}},  8'h80};
                    229 : data_out = {data_in[1087:864],  3'h7,  data_in[863:859],   8'h3,  {840{1'b0}},  8'h80};
                    230 : data_out = {data_in[1087:864],  2'h3,  data_in[863:858],   8'h7,  {840{1'b0}},  8'h80};
                    231 : data_out = {data_in[1087:864],  1'h1,  data_in[863:857],   8'hf,  {840{1'b0}},  8'h80};
                    232 : data_out = {data_in[1087:856],                             8'h1f, {840{1'b0}},  8'h80};

                    233 : data_out = {data_in[1087:856],  7'h1f, data_in[855],              {840{1'b0}},  8'h80};
                    234 : data_out = {data_in[1087:856],  6'h1f, data_in[855:854],          {840{1'b0}},  8'h80};
                    235 : data_out = {data_in[1087:856],  5'h1f, data_in[855:853],          {840{1'b0}},  8'h80};
                    236 : data_out = {data_in[1087:856],  4'hf,  data_in[855:852],   8'h1,  {832{1'b0}},  8'h80};
                    237 : data_out = {data_in[1087:856],  3'h7,  data_in[855:851],   8'h3,  {832{1'b0}},  8'h80};
                    238 : data_out = {data_in[1087:856],  2'h3,  data_in[855:850],   8'h7,  {832{1'b0}},  8'h80};
                    239 : data_out = {data_in[1087:856],  1'h1,  data_in[855:849],   8'hf,  {832{1'b0}},  8'h80};
                    240 : data_out = {data_in[1087:848],                             8'h1f, {832{1'b0}},  8'h80};

                    241 : data_out = {data_in[1087:848],  7'h1f, data_in[847],              {832{1'b0}},  8'h80};
                    242 : data_out = {data_in[1087:848],  6'h1f, data_in[847:846],          {832{1'b0}},  8'h80};
                    243 : data_out = {data_in[1087:848],  5'h1f, data_in[847:845],          {832{1'b0}},  8'h80};
                    244 : data_out = {data_in[1087:848],  4'hf,  data_in[847:844],   8'h1,  {824{1'b0}},  8'h80};
                    245 : data_out = {data_in[1087:848],  3'h7,  data_in[847:843],   8'h3,  {824{1'b0}},  8'h80};
                    246 : data_out = {data_in[1087:848],  2'h3,  data_in[847:842],   8'h7,  {824{1'b0}},  8'h80};
                    247 : data_out = {data_in[1087:848],  1'h1,  data_in[847:841],   8'hf,  {824{1'b0}},  8'h80};
                    248 : data_out = {data_in[1087:840],                             8'h1f, {824{1'b0}},  8'h80};

                    249 : data_out = {data_in[1087:840],  7'h1f, data_in[839],              {824{1'b0}},  8'h80};
                    250 : data_out = {data_in[1087:840],  6'h1f, data_in[839:838],          {824{1'b0}},  8'h80};
                    251 : data_out = {data_in[1087:840],  5'h1f, data_in[839:837],          {824{1'b0}},  8'h80};
                    252 : data_out = {data_in[1087:840],  4'hf,  data_in[839:836],   8'h1,  {816{1'b0}},  8'h80};
                    253 : data_out = {data_in[1087:840],  3'h7,  data_in[839:835],   8'h3,  {816{1'b0}},  8'h80};
                    254 : data_out = {data_in[1087:840],  2'h3,  data_in[839:834],   8'h7,  {816{1'b0}},  8'h80};
                    255 : data_out = {data_in[1087:840],  1'h1,  data_in[839:833],   8'hf,  {816{1'b0}},  8'h80};
                    256 : data_out = {data_in[1087:832],                             8'h1f, {816{1'b0}},  8'h80};

                    257 : data_out = {data_in[1087:832],  7'h1f, data_in[831],              {816{1'b0}},  8'h80};
                    258 : data_out = {data_in[1087:832],  6'h1f, data_in[831:830],          {816{1'b0}},  8'h80};
                    259 : data_out = {data_in[1087:832],  5'h1f, data_in[831:829],          {816{1'b0}},  8'h80};
                    260 : data_out = {data_in[1087:832],  4'hf,  data_in[831:828],   8'h1,  {808{1'b0}},  8'h80};
                    261 : data_out = {data_in[1087:832],  3'h7,  data_in[831:827],   8'h3,  {808{1'b0}},  8'h80};
                    262 : data_out = {data_in[1087:832],  2'h3,  data_in[831:826],   8'h7,  {808{1'b0}},  8'h80};
                    263 : data_out = {data_in[1087:832],  1'h1,  data_in[831:825],   8'hf,  {808{1'b0}},  8'h80};
                    264 : data_out = {data_in[1087:824],                             8'h1f, {808{1'b0}},  8'h80};

                    265 : data_out = {data_in[1087:824],  7'h1f, data_in[823],              {808{1'b0}},  8'h80};
                    266 : data_out = {data_in[1087:824],  6'h1f, data_in[823:822],          {808{1'b0}},  8'h80};
                    267 : data_out = {data_in[1087:824],  5'h1f, data_in[823:821],          {808{1'b0}},  8'h80};
                    268 : data_out = {data_in[1087:824],  4'hf,  data_in[823:820],   8'h1,  {800{1'b0}},  8'h80};
                    269 : data_out = {data_in[1087:824],  3'h7,  data_in[823:819],   8'h3,  {800{1'b0}},  8'h80};
                    270 : data_out = {data_in[1087:824],  2'h3,  data_in[823:818],   8'h7,  {800{1'b0}},  8'h80};
                    271 : data_out = {data_in[1087:824],  1'h1,  data_in[823:817],   8'hf,  {800{1'b0}},  8'h80};
                    272 : data_out = {data_in[1087:816],                             8'h1f, {800{1'b0}},  8'h80};

                    273 : data_out = {data_in[1087:816],  7'h1f, data_in[815],              {800{1'b0}},  8'h80};
                    274 : data_out = {data_in[1087:816],  6'h1f, data_in[815:814],          {800{1'b0}},  8'h80};
                    275 : data_out = {data_in[1087:816],  5'h1f, data_in[815:813],          {800{1'b0}},  8'h80};
                    276 : data_out = {data_in[1087:816],  4'hf,  data_in[815:812],   8'h1,  {792{1'b0}},  8'h80};
                    277 : data_out = {data_in[1087:816],  3'h7,  data_in[815:811],   8'h3,  {792{1'b0}},  8'h80};
                    278 : data_out = {data_in[1087:816],  2'h3,  data_in[815:810],   8'h7,  {792{1'b0}},  8'h80};
                    279 : data_out = {data_in[1087:816],  1'h1,  data_in[815:809],   8'hf,  {792{1'b0}},  8'h80};
                    280 : data_out = {data_in[1087:808],                             8'h1f, {792{1'b0}},  8'h80};

                    281 : data_out = {data_in[1087:808],  7'h1f, data_in[807],              {792{1'b0}},  8'h80};
                    282 : data_out = {data_in[1087:808],  6'h1f, data_in[807:806],          {792{1'b0}},  8'h80};
                    283 : data_out = {data_in[1087:808],  5'h1f, data_in[807:805],          {792{1'b0}},  8'h80};
                    284 : data_out = {data_in[1087:808],  4'hf,  data_in[807:804],   8'h1,  {784{1'b0}},  8'h80};
                    285 : data_out = {data_in[1087:808],  3'h7,  data_in[807:803],   8'h3,  {784{1'b0}},  8'h80};
                    286 : data_out = {data_in[1087:808],  2'h3,  data_in[807:802],   8'h7,  {784{1'b0}},  8'h80};
                    287 : data_out = {data_in[1087:808],  1'h1,  data_in[807:801],   8'hf,  {784{1'b0}},  8'h80};
                    288 : data_out = {data_in[1087:800],                             8'h1f, {784{1'b0}},  8'h80};

                    289 : data_out = {data_in[1087:800],  7'h1f, data_in[799],              {784{1'b0}},  8'h80};
                    290 : data_out = {data_in[1087:800],  6'h1f, data_in[799:798],          {784{1'b0}},  8'h80};
                    291 : data_out = {data_in[1087:800],  5'h1f, data_in[799:797],          {784{1'b0}},  8'h80};
                    292 : data_out = {data_in[1087:800],  4'hf,  data_in[799:796],   8'h1,  {776{1'b0}},  8'h80};
                    293 : data_out = {data_in[1087:800],  3'h7,  data_in[799:795],   8'h3,  {776{1'b0}},  8'h80};
                    294 : data_out = {data_in[1087:800],  2'h3,  data_in[799:794],   8'h7,  {776{1'b0}},  8'h80};
                    295 : data_out = {data_in[1087:800],  1'h1,  data_in[799:793],   8'hf,  {776{1'b0}},  8'h80};
                    296 : data_out = {data_in[1087:792],                             8'h1f, {776{1'b0}},  8'h80};

                    297 : data_out = {data_in[1087:792],  7'h1f, data_in[791],              {776{1'b0}},  8'h80};
                    298 : data_out = {data_in[1087:792],  6'h1f, data_in[791:790],          {776{1'b0}},  8'h80};
                    299 : data_out = {data_in[1087:792],  5'h1f, data_in[791:789],          {776{1'b0}},  8'h80};
                    300 : data_out = {data_in[1087:792],  4'hf,  data_in[791:788],   8'h1,  {768{1'b0}},  8'h80};
                    301 : data_out = {data_in[1087:792],  3'h7,  data_in[791:787],   8'h3,  {768{1'b0}},  8'h80};
                    302 : data_out = {data_in[1087:792],  2'h3,  data_in[791:786],   8'h7,  {768{1'b0}},  8'h80};
                    303 : data_out = {data_in[1087:792],  1'h1,  data_in[791:785],   8'hf,  {768{1'b0}},  8'h80};
                    304 : data_out = {data_in[1087:784],                             8'h1f, {768{1'b0}},  8'h80};

                    305 : data_out = {data_in[1087:784],  7'h1f, data_in[783],              {768{1'b0}},  8'h80};
                    306 : data_out = {data_in[1087:784],  6'h1f, data_in[783:782],          {768{1'b0}},  8'h80};
                    307 : data_out = {data_in[1087:784],  5'h1f, data_in[783:781],          {768{1'b0}},  8'h80};
                    308 : data_out = {data_in[1087:784],  4'hf,  data_in[783:780],   8'h1,  {760{1'b0}},  8'h80};
                    309 : data_out = {data_in[1087:784],  3'h7,  data_in[783:779],   8'h3,  {760{1'b0}},  8'h80};
                    310 : data_out = {data_in[1087:784],  2'h3,  data_in[783:778],   8'h7,  {760{1'b0}},  8'h80};
                    311 : data_out = {data_in[1087:784],  1'h1,  data_in[783:777],   8'hf,  {760{1'b0}},  8'h80};
                    312 : data_out = {data_in[1087:776],                             8'h1f, {760{1'b0}},  8'h80};

                    313 : data_out = {data_in[1087:776],  7'h1f, data_in[775],              {760{1'b0}},  8'h80};
                    314 : data_out = {data_in[1087:776],  6'h1f, data_in[775:774],          {760{1'b0}},  8'h80};
                    315 : data_out = {data_in[1087:776],  5'h1f, data_in[775:773],          {760{1'b0}},  8'h80};
                    316 : data_out = {data_in[1087:776],  4'hf,  data_in[775:772],   8'h1,  {752{1'b0}},  8'h80};
                    317 : data_out = {data_in[1087:776],  3'h7,  data_in[775:771],   8'h3,  {752{1'b0}},  8'h80};
                    318 : data_out = {data_in[1087:776],  2'h3,  data_in[775:770],   8'h7,  {752{1'b0}},  8'h80};
                    319 : data_out = {data_in[1087:776],  1'h1,  data_in[775:769],   8'hf,  {752{1'b0}},  8'h80};
                    320 : data_out = {data_in[1087:768],                             8'h1f, {752{1'b0}},  8'h80};

                    321 : data_out = {data_in[1087:768],  7'h1f, data_in[767],              {752{1'b0}},  8'h80};
                    322 : data_out = {data_in[1087:768],  6'h1f, data_in[767:766],          {752{1'b0}},  8'h80};
                    323 : data_out = {data_in[1087:768],  5'h1f, data_in[767:765],          {752{1'b0}},  8'h80};
                    324 : data_out = {data_in[1087:768],  4'hf,  data_in[767:764],   8'h1,  {744{1'b0}},  8'h80};
                    325 : data_out = {data_in[1087:768],  3'h7,  data_in[767:763],   8'h3,  {744{1'b0}},  8'h80};
                    326 : data_out = {data_in[1087:768],  2'h3,  data_in[767:762],   8'h7,  {744{1'b0}},  8'h80};
                    327 : data_out = {data_in[1087:768],  1'h1,  data_in[767:761],   8'hf,  {744{1'b0}},  8'h80};
                    328 : data_out = {data_in[1087:760],                             8'h1f, {744{1'b0}},  8'h80};

                    329 : data_out = {data_in[1087:760],  7'h1f, data_in[759],              {744{1'b0}},  8'h80};
                    330 : data_out = {data_in[1087:760],  6'h1f, data_in[759:758],          {744{1'b0}},  8'h80};
                    331 : data_out = {data_in[1087:760],  5'h1f, data_in[759:757],          {744{1'b0}},  8'h80};
                    332 : data_out = {data_in[1087:760],  4'hf,  data_in[759:756],   8'h1,  {736{1'b0}},  8'h80};
                    333 : data_out = {data_in[1087:760],  3'h7,  data_in[759:755],   8'h3,  {736{1'b0}},  8'h80};
                    334 : data_out = {data_in[1087:760],  2'h3,  data_in[759:754],   8'h7,  {736{1'b0}},  8'h80};
                    335 : data_out = {data_in[1087:760],  1'h1,  data_in[759:753],   8'hf,  {736{1'b0}},  8'h80};
                    336 : data_out = {data_in[1087:752],                             8'h1f, {736{1'b0}},  8'h80};

                    337 : data_out = {data_in[1087:752],  7'h1f, data_in[751],              {736{1'b0}},  8'h80};
                    338 : data_out = {data_in[1087:752],  6'h1f, data_in[751:750],          {736{1'b0}},  8'h80};
                    339 : data_out = {data_in[1087:752],  5'h1f, data_in[751:749],          {736{1'b0}},  8'h80};
                    340 : data_out = {data_in[1087:752],  4'hf,  data_in[751:748],   8'h1,  {728{1'b0}},  8'h80};
                    341 : data_out = {data_in[1087:752],  3'h7,  data_in[751:747],   8'h3,  {728{1'b0}},  8'h80};
                    342 : data_out = {data_in[1087:752],  2'h3,  data_in[751:746],   8'h7,  {728{1'b0}},  8'h80};
                    343 : data_out = {data_in[1087:752],  1'h1,  data_in[751:745],   8'hf,  {728{1'b0}},  8'h80};
                    344 : data_out = {data_in[1087:744],                             8'h1f, {728{1'b0}},  8'h80};

                    345 : data_out = {data_in[1087:744],  7'h1f, data_in[743],              {728{1'b0}},  8'h80};
                    346 : data_out = {data_in[1087:744],  6'h1f, data_in[743:742],          {728{1'b0}},  8'h80};
                    347 : data_out = {data_in[1087:744],  5'h1f, data_in[743:741],          {728{1'b0}},  8'h80};
                    348 : data_out = {data_in[1087:744],  4'hf,  data_in[743:740],   8'h1,  {720{1'b0}},  8'h80};
                    349 : data_out = {data_in[1087:744],  3'h7,  data_in[743:739],   8'h3,  {720{1'b0}},  8'h80};
                    350 : data_out = {data_in[1087:744],  2'h3,  data_in[743:738],   8'h7,  {720{1'b0}},  8'h80};
                    351 : data_out = {data_in[1087:744],  1'h1,  data_in[743:737],   8'hf,  {720{1'b0}},  8'h80};
                    352 : data_out = {data_in[1087:736],                             8'h1f, {720{1'b0}},  8'h80};

                    353 : data_out = {data_in[1087:736],  7'h1f, data_in[735],              {720{1'b0}},  8'h80};
                    354 : data_out = {data_in[1087:736],  6'h1f, data_in[735:734],          {720{1'b0}},  8'h80};
                    355 : data_out = {data_in[1087:736],  5'h1f, data_in[735:733],          {720{1'b0}},  8'h80};
                    356 : data_out = {data_in[1087:736],  4'hf,  data_in[735:732],   8'h1,  {712{1'b0}},  8'h80};
                    357 : data_out = {data_in[1087:736],  3'h7,  data_in[735:731],   8'h3,  {712{1'b0}},  8'h80};
                    358 : data_out = {data_in[1087:736],  2'h3,  data_in[735:730],   8'h7,  {712{1'b0}},  8'h80};
                    359 : data_out = {data_in[1087:736],  1'h1,  data_in[735:729],   8'hf,  {712{1'b0}},  8'h80};
                    360 : data_out = {data_in[1087:728],                             8'h1f, {712{1'b0}},  8'h80};

                    361 : data_out = {data_in[1087:728],  7'h1f, data_in[727],              {712{1'b0}},  8'h80};
                    362 : data_out = {data_in[1087:728],  6'h1f, data_in[727:726],          {712{1'b0}},  8'h80};
                    363 : data_out = {data_in[1087:728],  5'h1f, data_in[727:725],          {712{1'b0}},  8'h80};
                    364 : data_out = {data_in[1087:728],  4'hf,  data_in[727:724],   8'h1,  {704{1'b0}},  8'h80};
                    365 : data_out = {data_in[1087:728],  3'h7,  data_in[727:723],   8'h3,  {704{1'b0}},  8'h80};
                    366 : data_out = {data_in[1087:728],  2'h3,  data_in[727:722],   8'h7,  {704{1'b0}},  8'h80};
                    367 : data_out = {data_in[1087:728],  1'h1,  data_in[727:721],   8'hf,  {704{1'b0}},  8'h80};
                    368 : data_out = {data_in[1087:720],                             8'h1f, {704{1'b0}},  8'h80};

                    369 : data_out = {data_in[1087:720],  7'h1f, data_in[719],              {704{1'b0}},  8'h80};
                    370 : data_out = {data_in[1087:720],  6'h1f, data_in[719:718],          {704{1'b0}},  8'h80};
                    371 : data_out = {data_in[1087:720],  5'h1f, data_in[719:717],          {704{1'b0}},  8'h80};
                    372 : data_out = {data_in[1087:720],  4'hf,  data_in[719:716],   8'h1,  {696{1'b0}},  8'h80};
                    373 : data_out = {data_in[1087:720],  3'h7,  data_in[719:715],   8'h3,  {696{1'b0}},  8'h80};
                    374 : data_out = {data_in[1087:720],  2'h3,  data_in[719:714],   8'h7,  {696{1'b0}},  8'h80};
                    375 : data_out = {data_in[1087:720],  1'h1,  data_in[719:713],   8'hf,  {696{1'b0}},  8'h80};
                    376 : data_out = {data_in[1087:712],                             8'h1f, {696{1'b0}},  8'h80};

                    377 : data_out = {data_in[1087:712],  7'h1f, data_in[711],              {696{1'b0}},  8'h80};
                    378 : data_out = {data_in[1087:712],  6'h1f, data_in[711:710],          {696{1'b0}},  8'h80};
                    379 : data_out = {data_in[1087:712],  5'h1f, data_in[711:709],          {696{1'b0}},  8'h80};
                    380 : data_out = {data_in[1087:712],  4'hf,  data_in[711:708],   8'h1,  {688{1'b0}},  8'h80};
                    381 : data_out = {data_in[1087:712],  3'h7,  data_in[711:707],   8'h3,  {688{1'b0}},  8'h80};
                    382 : data_out = {data_in[1087:712],  2'h3,  data_in[711:706],   8'h7,  {688{1'b0}},  8'h80};
                    383 : data_out = {data_in[1087:712],  1'h1,  data_in[711:705],   8'hf,  {688{1'b0}},  8'h80};
                    384 : data_out = {data_in[1087:704],                             8'h1f, {688{1'b0}},  8'h80};

                    385 : data_out = {data_in[1087:704],  7'h1f, data_in[703],              {688{1'b0}},  8'h80};
                    386 : data_out = {data_in[1087:704],  6'h1f, data_in[703:702],          {688{1'b0}},  8'h80};
                    387 : data_out = {data_in[1087:704],  5'h1f, data_in[703:701],          {688{1'b0}},  8'h80};
                    388 : data_out = {data_in[1087:704],  4'hf,  data_in[703:700],   8'h1,  {680{1'b0}},  8'h80};
                    389 : data_out = {data_in[1087:704],  3'h7,  data_in[703:699],   8'h3,  {680{1'b0}},  8'h80};
                    390 : data_out = {data_in[1087:704],  2'h3,  data_in[703:698],   8'h7,  {680{1'b0}},  8'h80};
                    391 : data_out = {data_in[1087:704],  1'h1,  data_in[703:697],   8'hf,  {680{1'b0}},  8'h80};
                    392 : data_out = {data_in[1087:696],                             8'h1f, {680{1'b0}},  8'h80};

                    393 : data_out = {data_in[1087:696],  7'h1f, data_in[695],              {680{1'b0}},  8'h80};
                    394 : data_out = {data_in[1087:696],  6'h1f, data_in[695:694],          {680{1'b0}},  8'h80};
                    395 : data_out = {data_in[1087:696],  5'h1f, data_in[695:693],          {680{1'b0}},  8'h80};
                    396 : data_out = {data_in[1087:696],  4'hf,  data_in[695:692],   8'h1,  {672{1'b0}},  8'h80};
                    397 : data_out = {data_in[1087:696],  3'h7,  data_in[695:691],   8'h3,  {672{1'b0}},  8'h80};
                    398 : data_out = {data_in[1087:696],  2'h3,  data_in[695:690],   8'h7,  {672{1'b0}},  8'h80};
                    399 : data_out = {data_in[1087:696],  1'h1,  data_in[695:689],   8'hf,  {672{1'b0}},  8'h80};
                    400 : data_out = {data_in[1087:688],                             8'h1f, {672{1'b0}},  8'h80};

                    401 : data_out = {data_in[1087:688],  7'h1f, data_in[687],              {672{1'b0}},  8'h80};
                    402 : data_out = {data_in[1087:688],  6'h1f, data_in[687:686],          {672{1'b0}},  8'h80};
                    403 : data_out = {data_in[1087:688],  5'h1f, data_in[687:685],          {672{1'b0}},  8'h80};
                    404 : data_out = {data_in[1087:688],  4'hf,  data_in[687:684],   8'h1,  {664{1'b0}},  8'h80};
                    405 : data_out = {data_in[1087:688],  3'h7,  data_in[687:683],   8'h3,  {664{1'b0}},  8'h80};
                    406 : data_out = {data_in[1087:688],  2'h3,  data_in[687:682],   8'h7,  {664{1'b0}},  8'h80};
                    407 : data_out = {data_in[1087:688],  1'h1,  data_in[687:681],   8'hf,  {664{1'b0}},  8'h80};
                    408 : data_out = {data_in[1087:680],                             8'h1f, {664{1'b0}},  8'h80};

                    409 : data_out = {data_in[1087:680],  7'h1f, data_in[679],              {664{1'b0}},  8'h80};
                    410 : data_out = {data_in[1087:680],  6'h1f, data_in[679:678],          {664{1'b0}},  8'h80};
                    411 : data_out = {data_in[1087:680],  5'h1f, data_in[679:677],          {664{1'b0}},  8'h80};
                    412 : data_out = {data_in[1087:680],  4'hf,  data_in[679:676],   8'h1,  {656{1'b0}},  8'h80};
                    413 : data_out = {data_in[1087:680],  3'h7,  data_in[679:675],   8'h3,  {656{1'b0}},  8'h80};
                    414 : data_out = {data_in[1087:680],  2'h3,  data_in[679:674],   8'h7,  {656{1'b0}},  8'h80};
                    415 : data_out = {data_in[1087:680],  1'h1,  data_in[679:673],   8'hf,  {656{1'b0}},  8'h80};
                    416 : data_out = {data_in[1087:672],                             8'h1f, {656{1'b0}},  8'h80};

                    417 : data_out = {data_in[1087:672],  7'h1f, data_in[671],              {656{1'b0}},  8'h80};
                    418 : data_out = {data_in[1087:672],  6'h1f, data_in[671:670],          {656{1'b0}},  8'h80};
                    419 : data_out = {data_in[1087:672],  5'h1f, data_in[671:669],          {656{1'b0}},  8'h80};
                    420 : data_out = {data_in[1087:672],  4'hf,  data_in[671:668],   8'h1,  {648{1'b0}},  8'h80};
                    421 : data_out = {data_in[1087:672],  3'h7,  data_in[671:667],   8'h3,  {648{1'b0}},  8'h80};
                    422 : data_out = {data_in[1087:672],  2'h3,  data_in[671:666],   8'h7,  {648{1'b0}},  8'h80};
                    423 : data_out = {data_in[1087:672],  1'h1,  data_in[671:665],   8'hf,  {648{1'b0}},  8'h80};
                    424 : data_out = {data_in[1087:664],                             8'h1f, {648{1'b0}},  8'h80};

                    425 : data_out = {data_in[1087:664],  7'h1f, data_in[663],              {648{1'b0}},  8'h80};
                    426 : data_out = {data_in[1087:664],  6'h1f, data_in[663:662],          {648{1'b0}},  8'h80};
                    427 : data_out = {data_in[1087:664],  5'h1f, data_in[663:661],          {648{1'b0}},  8'h80};
                    428 : data_out = {data_in[1087:664],  4'hf,  data_in[663:660],   8'h1,  {640{1'b0}},  8'h80};
                    429 : data_out = {data_in[1087:664],  3'h7,  data_in[663:659],   8'h3,  {640{1'b0}},  8'h80};
                    430 : data_out = {data_in[1087:664],  2'h3,  data_in[663:658],   8'h7,  {640{1'b0}},  8'h80};
                    431 : data_out = {data_in[1087:664],  1'h1,  data_in[663:657],   8'hf,  {640{1'b0}},  8'h80};
                    432 : data_out = {data_in[1087:656],                             8'h1f, {640{1'b0}},  8'h80};

                    433 : data_out = {data_in[1087:656],  7'h1f, data_in[655],              {640{1'b0}},  8'h80};
                    434 : data_out = {data_in[1087:656],  6'h1f, data_in[655:654],          {640{1'b0}},  8'h80};
                    435 : data_out = {data_in[1087:656],  5'h1f, data_in[655:653],          {640{1'b0}},  8'h80};
                    436 : data_out = {data_in[1087:656],  4'hf,  data_in[655:652],   8'h1,  {632{1'b0}},  8'h80};
                    437 : data_out = {data_in[1087:656],  3'h7,  data_in[655:651],   8'h3,  {632{1'b0}},  8'h80};
                    438 : data_out = {data_in[1087:656],  2'h3,  data_in[655:650],   8'h7,  {632{1'b0}},  8'h80};
                    439 : data_out = {data_in[1087:656],  1'h1,  data_in[655:649],   8'hf,  {632{1'b0}},  8'h80};
                    440 : data_out = {data_in[1087:648],                             8'h1f, {632{1'b0}},  8'h80};

                    441 : data_out = {data_in[1087:648],  7'h1f, data_in[647],              {632{1'b0}},  8'h80};
                    442 : data_out = {data_in[1087:648],  6'h1f, data_in[647:646],          {632{1'b0}},  8'h80};
                    443 : data_out = {data_in[1087:648],  5'h1f, data_in[647:645],          {632{1'b0}},  8'h80};
                    444 : data_out = {data_in[1087:648],  4'hf,  data_in[647:644],   8'h1,  {624{1'b0}},  8'h80};
                    445 : data_out = {data_in[1087:648],  3'h7,  data_in[647:643],   8'h3,  {624{1'b0}},  8'h80};
                    446 : data_out = {data_in[1087:648],  2'h3,  data_in[647:642],   8'h7,  {624{1'b0}},  8'h80};
                    447 : data_out = {data_in[1087:648],  1'h1,  data_in[647:641],   8'hf,  {624{1'b0}},  8'h80};
                    448 : data_out = {data_in[1087:640],                             8'h1f, {624{1'b0}},  8'h80};

                    449 : data_out = {data_in[1087:640],  7'h1f, data_in[639],              {624{1'b0}},  8'h80};
                    450 : data_out = {data_in[1087:640],  6'h1f, data_in[639:638],          {624{1'b0}},  8'h80};
                    451 : data_out = {data_in[1087:640],  5'h1f, data_in[639:637],          {624{1'b0}},  8'h80};
                    452 : data_out = {data_in[1087:640],  4'hf,  data_in[639:636],   8'h1,  {616{1'b0}},  8'h80};
                    453 : data_out = {data_in[1087:640],  3'h7,  data_in[639:635],   8'h3,  {616{1'b0}},  8'h80};
                    454 : data_out = {data_in[1087:640],  2'h3,  data_in[639:634],   8'h7,  {616{1'b0}},  8'h80};
                    455 : data_out = {data_in[1087:640],  1'h1,  data_in[639:633],   8'hf,  {616{1'b0}},  8'h80};
                    456 : data_out = {data_in[1087:632],                             8'h1f, {616{1'b0}},  8'h80};

                    457 : data_out = {data_in[1087:632],  7'h1f, data_in[631],              {616{1'b0}},  8'h80};
                    458 : data_out = {data_in[1087:632],  6'h1f, data_in[631:630],          {616{1'b0}},  8'h80};
                    459 : data_out = {data_in[1087:632],  5'h1f, data_in[631:629],          {616{1'b0}},  8'h80};
                    460 : data_out = {data_in[1087:632],  4'hf,  data_in[631:628],   8'h1,  {608{1'b0}},  8'h80};
                    461 : data_out = {data_in[1087:632],  3'h7,  data_in[631:627],   8'h3,  {608{1'b0}},  8'h80};
                    462 : data_out = {data_in[1087:632],  2'h3,  data_in[631:626],   8'h7,  {608{1'b0}},  8'h80};
                    463 : data_out = {data_in[1087:632],  1'h1,  data_in[631:625],   8'hf,  {608{1'b0}},  8'h80};
                    464 : data_out = {data_in[1087:624],                             8'h1f, {608{1'b0}},  8'h80};

                    465 : data_out = {data_in[1087:624],  7'h1f, data_in[623],              {608{1'b0}},  8'h80};
                    466 : data_out = {data_in[1087:624],  6'h1f, data_in[623:622],          {608{1'b0}},  8'h80};
                    467 : data_out = {data_in[1087:624],  5'h1f, data_in[623:621],          {608{1'b0}},  8'h80};
                    468 : data_out = {data_in[1087:624],  4'hf,  data_in[623:620],   8'h1,  {600{1'b0}},  8'h80};
                    469 : data_out = {data_in[1087:624],  3'h7,  data_in[623:619],   8'h3,  {600{1'b0}},  8'h80};
                    470 : data_out = {data_in[1087:624],  2'h3,  data_in[623:618],   8'h7,  {600{1'b0}},  8'h80};
                    471 : data_out = {data_in[1087:624],  1'h1,  data_in[623:617],   8'hf,  {600{1'b0}},  8'h80};
                    472 : data_out = {data_in[1087:616],                             8'h1f, {600{1'b0}},  8'h80};

                    473 : data_out = {data_in[1087:616],  7'h1f, data_in[615],              {600{1'b0}},  8'h80};
                    474 : data_out = {data_in[1087:616],  6'h1f, data_in[615:614],          {600{1'b0}},  8'h80};
                    475 : data_out = {data_in[1087:616],  5'h1f, data_in[615:613],          {600{1'b0}},  8'h80};
                    476 : data_out = {data_in[1087:616],  4'hf,  data_in[615:612],   8'h1,  {592{1'b0}},  8'h80};
                    477 : data_out = {data_in[1087:616],  3'h7,  data_in[615:611],   8'h3,  {592{1'b0}},  8'h80};
                    478 : data_out = {data_in[1087:616],  2'h3,  data_in[615:610],   8'h7,  {592{1'b0}},  8'h80};
                    479 : data_out = {data_in[1087:616],  1'h1,  data_in[615:609],   8'hf,  {592{1'b0}},  8'h80};
                    480 : data_out = {data_in[1087:608],                             8'h1f, {592{1'b0}},  8'h80};

                    481 : data_out = {data_in[1087:608],  7'h1f, data_in[607],              {592{1'b0}},  8'h80};
                    482 : data_out = {data_in[1087:608],  6'h1f, data_in[607:606],          {592{1'b0}},  8'h80};
                    483 : data_out = {data_in[1087:608],  5'h1f, data_in[607:605],          {592{1'b0}},  8'h80};
                    484 : data_out = {data_in[1087:608],  4'hf,  data_in[607:604],   8'h1,  {584{1'b0}},  8'h80};
                    485 : data_out = {data_in[1087:608],  3'h7,  data_in[607:603],   8'h3,  {584{1'b0}},  8'h80};
                    486 : data_out = {data_in[1087:608],  2'h3,  data_in[607:602],   8'h7,  {584{1'b0}},  8'h80};
                    487 : data_out = {data_in[1087:608],  1'h1,  data_in[607:601],   8'hf,  {584{1'b0}},  8'h80};
                    488 : data_out = {data_in[1087:600],                             8'h1f, {584{1'b0}},  8'h80};

                    489 : data_out = {data_in[1087:600],  7'h1f, data_in[599],              {584{1'b0}},  8'h80};
                    490 : data_out = {data_in[1087:600],  6'h1f, data_in[599:598],          {584{1'b0}},  8'h80};
                    491 : data_out = {data_in[1087:600],  5'h1f, data_in[599:597],          {584{1'b0}},  8'h80};
                    492 : data_out = {data_in[1087:600],  4'hf,  data_in[599:596],   8'h1,  {576{1'b0}},  8'h80};
                    493 : data_out = {data_in[1087:600],  3'h7,  data_in[599:595],   8'h3,  {576{1'b0}},  8'h80};
                    494 : data_out = {data_in[1087:600],  2'h3,  data_in[599:594],   8'h7,  {576{1'b0}},  8'h80};
                    495 : data_out = {data_in[1087:600],  1'h1,  data_in[599:593],   8'hf,  {576{1'b0}},  8'h80};
                    496 : data_out = {data_in[1087:592],                             8'h1f, {576{1'b0}},  8'h80};

                    497 : data_out = {data_in[1087:592],  7'h1f, data_in[591],              {576{1'b0}},  8'h80};
                    498 : data_out = {data_in[1087:592],  6'h1f, data_in[591:590],          {576{1'b0}},  8'h80};
                    499 : data_out = {data_in[1087:592],  5'h1f, data_in[591:589],          {576{1'b0}},  8'h80};
                    500 : data_out = {data_in[1087:592],  4'hf,  data_in[591:588],   8'h1,  {568{1'b0}},  8'h80};
                    501 : data_out = {data_in[1087:592],  3'h7,  data_in[591:587],   8'h3,  {568{1'b0}},  8'h80};
                    502 : data_out = {data_in[1087:592],  2'h3,  data_in[591:586],   8'h7,  {568{1'b0}},  8'h80};
                    503 : data_out = {data_in[1087:592],  1'h1,  data_in[591:585],   8'hf,  {568{1'b0}},  8'h80};
                    504 : data_out = {data_in[1087:584],                             8'h1f, {568{1'b0}},  8'h80};

                    505 : data_out = {data_in[1087:584],  7'h1f, data_in[583],              {568{1'b0}},  8'h80};
                    506 : data_out = {data_in[1087:584],  6'h1f, data_in[583:582],          {568{1'b0}},  8'h80};
                    507 : data_out = {data_in[1087:584],  5'h1f, data_in[583:581],          {568{1'b0}},  8'h80};
                    508 : data_out = {data_in[1087:584],  4'hf,  data_in[583:580],   8'h1,  {560{1'b0}},  8'h80};
                    509 : data_out = {data_in[1087:584],  3'h7,  data_in[583:579],   8'h3,  {560{1'b0}},  8'h80};
                    510 : data_out = {data_in[1087:584],  2'h3,  data_in[583:578],   8'h7,  {560{1'b0}},  8'h80};
                    511 : data_out = {data_in[1087:584],  1'h1,  data_in[583:577],   8'hf,  {560{1'b0}},  8'h80};
                    512 : data_out = {data_in[1087:576],                             8'h1f, {560{1'b0}},  8'h80};

                    513 : data_out = {data_in[1087:576],  7'h1f, data_in[575],              {560{1'b0}},  8'h80};
                    514 : data_out = {data_in[1087:576],  6'h1f, data_in[575:574],          {560{1'b0}},  8'h80};
                    515 : data_out = {data_in[1087:576],  5'h1f, data_in[575:573],          {560{1'b0}},  8'h80};
                    516 : data_out = {data_in[1087:576],  4'hf,  data_in[575:572],   8'h1,  {552{1'b0}},  8'h80};
                    517 : data_out = {data_in[1087:576],  3'h7,  data_in[575:571],   8'h3,  {552{1'b0}},  8'h80};
                    518 : data_out = {data_in[1087:576],  2'h3,  data_in[575:570],   8'h7,  {552{1'b0}},  8'h80};
                    519 : data_out = {data_in[1087:576],  1'h1,  data_in[575:569],   8'hf,  {552{1'b0}},  8'h80};
                    520 : data_out = {data_in[1087:568],                             8'h1f, {552{1'b0}},  8'h80};

                    521 : data_out = {data_in[1087:568],  7'h1f, data_in[567],              {552{1'b0}},  8'h80};
                    522 : data_out = {data_in[1087:568],  6'h1f, data_in[567:566],          {552{1'b0}},  8'h80};
                    523 : data_out = {data_in[1087:568],  5'h1f, data_in[567:565],          {552{1'b0}},  8'h80};
                    524 : data_out = {data_in[1087:568],  4'hf,  data_in[567:564],   8'h1,  {544{1'b0}},  8'h80};
                    525 : data_out = {data_in[1087:568],  3'h7,  data_in[567:563],   8'h3,  {544{1'b0}},  8'h80};
                    526 : data_out = {data_in[1087:568],  2'h3,  data_in[567:562],   8'h7,  {544{1'b0}},  8'h80};
                    527 : data_out = {data_in[1087:568],  1'h1,  data_in[567:561],   8'hf,  {544{1'b0}},  8'h80};
                    528 : data_out = {data_in[1087:560],                             8'h1f, {544{1'b0}},  8'h80};

                    529 : data_out = {data_in[1087:560],  7'h1f, data_in[559],              {544{1'b0}},  8'h80};
                    530 : data_out = {data_in[1087:560],  6'h1f, data_in[559:558],          {544{1'b0}},  8'h80};
                    531 : data_out = {data_in[1087:560],  5'h1f, data_in[559:557],          {544{1'b0}},  8'h80};
                    532 : data_out = {data_in[1087:560],  4'hf,  data_in[559:556],   8'h1,  {536{1'b0}},  8'h80};
                    533 : data_out = {data_in[1087:560],  3'h7,  data_in[559:555],   8'h3,  {536{1'b0}},  8'h80};
                    534 : data_out = {data_in[1087:560],  2'h3,  data_in[559:554],   8'h7,  {536{1'b0}},  8'h80};
                    535 : data_out = {data_in[1087:560],  1'h1,  data_in[559:553],   8'hf,  {536{1'b0}},  8'h80};
                    536 : data_out = {data_in[1087:552],                             8'h1f, {536{1'b0}},  8'h80};

                    537 : data_out = {data_in[1087:552],  7'h1f, data_in[551],              {536{1'b0}},  8'h80};
                    538 : data_out = {data_in[1087:552],  6'h1f, data_in[551:550],          {536{1'b0}},  8'h80};
                    539 : data_out = {data_in[1087:552],  5'h1f, data_in[551:549],          {536{1'b0}},  8'h80};
                    540 : data_out = {data_in[1087:552],  4'hf,  data_in[551:548],   8'h1,  {528{1'b0}},  8'h80};
                    541 : data_out = {data_in[1087:552],  3'h7,  data_in[551:547],   8'h3,  {528{1'b0}},  8'h80};
                    542 : data_out = {data_in[1087:552],  2'h3,  data_in[551:546],   8'h7,  {528{1'b0}},  8'h80};
                    543 : data_out = {data_in[1087:552],  1'h1,  data_in[551:545],   8'hf,  {528{1'b0}},  8'h80};
                    544 : data_out = {data_in[1087:544],                             8'h1f, {528{1'b0}},  8'h80};

                    545 : data_out = {data_in[1087:544],  7'h1f, data_in[543],              {528{1'b0}},  8'h80};
                    546 : data_out = {data_in[1087:544],  6'h1f, data_in[543:542],          {528{1'b0}},  8'h80};
                    547 : data_out = {data_in[1087:544],  5'h1f, data_in[543:541],          {528{1'b0}},  8'h80};
                    548 : data_out = {data_in[1087:544],  4'hf,  data_in[543:540],   8'h1,  {520{1'b0}},  8'h80};
                    549 : data_out = {data_in[1087:544],  3'h7,  data_in[543:539],   8'h3,  {520{1'b0}},  8'h80};
                    550 : data_out = {data_in[1087:544],  2'h3,  data_in[543:538],   8'h7,  {520{1'b0}},  8'h80};
                    551 : data_out = {data_in[1087:544],  1'h1,  data_in[543:537],   8'hf,  {520{1'b0}},  8'h80};
                    552 : data_out = {data_in[1087:536],                             8'h1f, {520{1'b0}},  8'h80};

                    553 : data_out = {data_in[1087:536],  7'h1f, data_in[535],              {520{1'b0}},  8'h80};
                    554 : data_out = {data_in[1087:536],  6'h1f, data_in[535:534],          {520{1'b0}},  8'h80};
                    555 : data_out = {data_in[1087:536],  5'h1f, data_in[535:533],          {520{1'b0}},  8'h80};
                    556 : data_out = {data_in[1087:536],  4'hf,  data_in[535:532],   8'h1,  {512{1'b0}},  8'h80};
                    557 : data_out = {data_in[1087:536],  3'h7,  data_in[535:531],   8'h3,  {512{1'b0}},  8'h80};
                    558 : data_out = {data_in[1087:536],  2'h3,  data_in[535:530],   8'h7,  {512{1'b0}},  8'h80};
                    559 : data_out = {data_in[1087:536],  1'h1,  data_in[535:529],   8'hf,  {512{1'b0}},  8'h80};
                    560 : data_out = {data_in[1087:528],                             8'h1f, {512{1'b0}},  8'h80};

                    561 : data_out = {data_in[1087:528],  7'h1f, data_in[527],              {512{1'b0}},  8'h80};
                    562 : data_out = {data_in[1087:528],  6'h1f, data_in[527:526],          {512{1'b0}},  8'h80};
                    563 : data_out = {data_in[1087:528],  5'h1f, data_in[527:525],          {512{1'b0}},  8'h80};
                    564 : data_out = {data_in[1087:528],  4'hf,  data_in[527:524],   8'h1,  {504{1'b0}},  8'h80};
                    565 : data_out = {data_in[1087:528],  3'h7,  data_in[527:523],   8'h3,  {504{1'b0}},  8'h80};
                    566 : data_out = {data_in[1087:528],  2'h3,  data_in[527:522],   8'h7,  {504{1'b0}},  8'h80};
                    567 : data_out = {data_in[1087:528],  1'h1,  data_in[527:521],   8'hf,  {504{1'b0}},  8'h80};
                    568 : data_out = {data_in[1087:520],                             8'h1f, {504{1'b0}},  8'h80};

                    569 : data_out = {data_in[1087:520],  7'h1f, data_in[519],              {504{1'b0}},  8'h80};
                    570 : data_out = {data_in[1087:520],  6'h1f, data_in[519:518],          {504{1'b0}},  8'h80};
                    571 : data_out = {data_in[1087:520],  5'h1f, data_in[519:517],          {504{1'b0}},  8'h80};
                    572 : data_out = {data_in[1087:520],  4'hf,  data_in[519:516],   8'h1,  {496{1'b0}},  8'h80};
                    573 : data_out = {data_in[1087:520],  3'h7,  data_in[519:515],   8'h3,  {496{1'b0}},  8'h80};
                    574 : data_out = {data_in[1087:520],  2'h3,  data_in[519:514],   8'h7,  {496{1'b0}},  8'h80};
                    575 : data_out = {data_in[1087:520],  1'h1,  data_in[519:513],   8'hf,  {496{1'b0}},  8'h80};
                    576 : data_out = {data_in[1087:512],                             8'h1f, {496{1'b0}},  8'h80};

                    577 : data_out = {data_in[1087:512],  7'h1f, data_in[511],              {496{1'b0}},  8'h80};
                    578 : data_out = {data_in[1087:512],  6'h1f, data_in[511:510],          {496{1'b0}},  8'h80};
                    579 : data_out = {data_in[1087:512],  5'h1f, data_in[511:509],          {496{1'b0}},  8'h80};
                    580 : data_out = {data_in[1087:512],  4'hf,  data_in[511:508],   8'h1,  {488{1'b0}},  8'h80};
                    581 : data_out = {data_in[1087:512],  3'h7,  data_in[511:507],   8'h3,  {488{1'b0}},  8'h80};
                    582 : data_out = {data_in[1087:512],  2'h3,  data_in[511:506],   8'h7,  {488{1'b0}},  8'h80};
                    583 : data_out = {data_in[1087:512],  1'h1,  data_in[511:505],   8'hf,  {488{1'b0}},  8'h80};
                    584 : data_out = {data_in[1087:504],                             8'h1f, {488{1'b0}},  8'h80};

                    585 : data_out = {data_in[1087:504],  7'h1f, data_in[503],              {488{1'b0}},  8'h80};
                    586 : data_out = {data_in[1087:504],  6'h1f, data_in[503:502],          {488{1'b0}},  8'h80};
                    587 : data_out = {data_in[1087:504],  5'h1f, data_in[503:501],          {488{1'b0}},  8'h80};
                    588 : data_out = {data_in[1087:504],  4'hf,  data_in[503:500],   8'h1,  {480{1'b0}},  8'h80};
                    589 : data_out = {data_in[1087:504],  3'h7,  data_in[503:499],   8'h3,  {480{1'b0}},  8'h80};
                    590 : data_out = {data_in[1087:504],  2'h3,  data_in[503:498],   8'h7,  {480{1'b0}},  8'h80};
                    591 : data_out = {data_in[1087:504],  1'h1,  data_in[503:497],   8'hf,  {480{1'b0}},  8'h80};
                    592 : data_out = {data_in[1087:496],                             8'h1f, {480{1'b0}},  8'h80};

                    593 : data_out = {data_in[1087:496],  7'h1f, data_in[495],              {480{1'b0}},  8'h80};
                    594 : data_out = {data_in[1087:496],  6'h1f, data_in[495:494],          {480{1'b0}},  8'h80};
                    595 : data_out = {data_in[1087:496],  5'h1f, data_in[495:493],          {480{1'b0}},  8'h80};
                    596 : data_out = {data_in[1087:496],  4'hf,  data_in[495:492],   8'h1,  {472{1'b0}},  8'h80};
                    597 : data_out = {data_in[1087:496],  3'h7,  data_in[495:491],   8'h3,  {472{1'b0}},  8'h80};
                    598 : data_out = {data_in[1087:496],  2'h3,  data_in[495:490],   8'h7,  {472{1'b0}},  8'h80};
                    599 : data_out = {data_in[1087:496],  1'h1,  data_in[495:489],   8'hf,  {472{1'b0}},  8'h80};
                    600 : data_out = {data_in[1087:488],                             8'h1f, {472{1'b0}},  8'h80};

                    601 : data_out = {data_in[1087:488],  7'h1f, data_in[487],              {472{1'b0}},  8'h80};
                    602 : data_out = {data_in[1087:488],  6'h1f, data_in[487:486],          {472{1'b0}},  8'h80};
                    603 : data_out = {data_in[1087:488],  5'h1f, data_in[487:485],          {472{1'b0}},  8'h80};
                    604 : data_out = {data_in[1087:488],  4'hf,  data_in[487:484],   8'h1,  {464{1'b0}},  8'h80};
                    605 : data_out = {data_in[1087:488],  3'h7,  data_in[487:483],   8'h3,  {464{1'b0}},  8'h80};
                    606 : data_out = {data_in[1087:488],  2'h3,  data_in[487:482],   8'h7,  {464{1'b0}},  8'h80};
                    607 : data_out = {data_in[1087:488],  1'h1,  data_in[487:481],   8'hf,  {464{1'b0}},  8'h80};
                    608 : data_out = {data_in[1087:480],                             8'h1f, {464{1'b0}},  8'h80};

                    609 : data_out = {data_in[1087:480],  7'h1f, data_in[479],              {464{1'b0}},  8'h80};
                    610 : data_out = {data_in[1087:480],  6'h1f, data_in[479:478],          {464{1'b0}},  8'h80};
                    611 : data_out = {data_in[1087:480],  5'h1f, data_in[479:477],          {464{1'b0}},  8'h80};
                    612 : data_out = {data_in[1087:480],  4'hf,  data_in[479:476],   8'h1,  {456{1'b0}},  8'h80};
                    613 : data_out = {data_in[1087:480],  3'h7,  data_in[479:475],   8'h3,  {456{1'b0}},  8'h80};
                    614 : data_out = {data_in[1087:480],  2'h3,  data_in[479:474],   8'h7,  {456{1'b0}},  8'h80};
                    615 : data_out = {data_in[1087:480],  1'h1,  data_in[479:473],   8'hf,  {456{1'b0}},  8'h80};
                    616 : data_out = {data_in[1087:472],                             8'h1f, {456{1'b0}},  8'h80};

                    617 : data_out = {data_in[1087:472],  7'h1f, data_in[471],              {456{1'b0}},  8'h80};
                    618 : data_out = {data_in[1087:472],  6'h1f, data_in[471:470],          {456{1'b0}},  8'h80};
                    619 : data_out = {data_in[1087:472],  5'h1f, data_in[471:469],          {456{1'b0}},  8'h80};
                    620 : data_out = {data_in[1087:472],  4'hf,  data_in[471:468],   8'h1,  {448{1'b0}},  8'h80};
                    621 : data_out = {data_in[1087:472],  3'h7,  data_in[471:467],   8'h3,  {448{1'b0}},  8'h80};
                    622 : data_out = {data_in[1087:472],  2'h3,  data_in[471:466],   8'h7,  {448{1'b0}},  8'h80};
                    623 : data_out = {data_in[1087:472],  1'h1,  data_in[471:465],   8'hf,  {448{1'b0}},  8'h80};
                    624 : data_out = {data_in[1087:464],                             8'h1f, {448{1'b0}},  8'h80};

                    625 : data_out = {data_in[1087:464],  7'h1f, data_in[463],              {448{1'b0}},  8'h80};
                    626 : data_out = {data_in[1087:464],  6'h1f, data_in[463:462],          {448{1'b0}},  8'h80};
                    627 : data_out = {data_in[1087:464],  5'h1f, data_in[463:461],          {448{1'b0}},  8'h80};
                    628 : data_out = {data_in[1087:464],  4'hf,  data_in[463:460],   8'h1,  {440{1'b0}},  8'h80};
                    629 : data_out = {data_in[1087:464],  3'h7,  data_in[463:459],   8'h3,  {440{1'b0}},  8'h80};
                    630 : data_out = {data_in[1087:464],  2'h3,  data_in[463:458],   8'h7,  {440{1'b0}},  8'h80};
                    631 : data_out = {data_in[1087:464],  1'h1,  data_in[463:457],   8'hf,  {440{1'b0}},  8'h80};
                    632 : data_out = {data_in[1087:456],                             8'h1f, {440{1'b0}},  8'h80};

                    633 : data_out = {data_in[1087:456],  7'h1f, data_in[455],              {440{1'b0}},  8'h80};
                    634 : data_out = {data_in[1087:456],  6'h1f, data_in[455:454],          {440{1'b0}},  8'h80};
                    635 : data_out = {data_in[1087:456],  5'h1f, data_in[455:453],          {440{1'b0}},  8'h80};
                    636 : data_out = {data_in[1087:456],  4'hf,  data_in[455:452],   8'h1,  {432{1'b0}},  8'h80};
                    637 : data_out = {data_in[1087:456],  3'h7,  data_in[455:451],   8'h3,  {432{1'b0}},  8'h80};
                    638 : data_out = {data_in[1087:456],  2'h3,  data_in[455:450],   8'h7,  {432{1'b0}},  8'h80};
                    639 : data_out = {data_in[1087:456],  1'h1,  data_in[455:449],   8'hf,  {432{1'b0}},  8'h80};
                    640 : data_out = {data_in[1087:448],                             8'h1f, {432{1'b0}},  8'h80};

                    641 : data_out = {data_in[1087:448],  7'h1f, data_in[447],              {432{1'b0}},  8'h80};
                    642 : data_out = {data_in[1087:448],  6'h1f, data_in[447:446],          {432{1'b0}},  8'h80};
                    643 : data_out = {data_in[1087:448],  5'h1f, data_in[447:445],          {432{1'b0}},  8'h80};
                    644 : data_out = {data_in[1087:448],  4'hf,  data_in[447:444],   8'h1,  {424{1'b0}},  8'h80};
                    645 : data_out = {data_in[1087:448],  3'h7,  data_in[447:443],   8'h3,  {424{1'b0}},  8'h80};
                    646 : data_out = {data_in[1087:448],  2'h3,  data_in[447:442],   8'h7,  {424{1'b0}},  8'h80};
                    647 : data_out = {data_in[1087:448],  1'h1,  data_in[447:441],   8'hf,  {424{1'b0}},  8'h80};
                    648 : data_out = {data_in[1087:440],                             8'h1f, {424{1'b0}},  8'h80};

                    649 : data_out = {data_in[1087:440],  7'h1f, data_in[439],              {424{1'b0}},  8'h80};
                    650 : data_out = {data_in[1087:440],  6'h1f, data_in[439:438],          {424{1'b0}},  8'h80};
                    651 : data_out = {data_in[1087:440],  5'h1f, data_in[439:437],          {424{1'b0}},  8'h80};
                    652 : data_out = {data_in[1087:440],  4'hf,  data_in[439:436],   8'h1,  {416{1'b0}},  8'h80};
                    653 : data_out = {data_in[1087:440],  3'h7,  data_in[439:435],   8'h3,  {416{1'b0}},  8'h80};
                    654 : data_out = {data_in[1087:440],  2'h3,  data_in[439:434],   8'h7,  {416{1'b0}},  8'h80};
                    655 : data_out = {data_in[1087:440],  1'h1,  data_in[439:433],   8'hf,  {416{1'b0}},  8'h80};
                    656 : data_out = {data_in[1087:432],                             8'h1f, {416{1'b0}},  8'h80};

                    657 : data_out = {data_in[1087:432],  7'h1f, data_in[431],              {416{1'b0}},  8'h80};
                    658 : data_out = {data_in[1087:432],  6'h1f, data_in[431:430],          {416{1'b0}},  8'h80};
                    659 : data_out = {data_in[1087:432],  5'h1f, data_in[431:429],          {416{1'b0}},  8'h80};
                    660 : data_out = {data_in[1087:432],  4'hf,  data_in[431:428],   8'h1,  {408{1'b0}},  8'h80};
                    661 : data_out = {data_in[1087:432],  3'h7,  data_in[431:427],   8'h3,  {408{1'b0}},  8'h80};
                    662 : data_out = {data_in[1087:432],  2'h3,  data_in[431:426],   8'h7,  {408{1'b0}},  8'h80};
                    663 : data_out = {data_in[1087:432],  1'h1,  data_in[431:425],   8'hf,  {408{1'b0}},  8'h80};
                    664 : data_out = {data_in[1087:424],                             8'h1f, {408{1'b0}},  8'h80};

                    665 : data_out = {data_in[1087:424],  7'h1f, data_in[423],              {408{1'b0}},  8'h80};
                    666 : data_out = {data_in[1087:424],  6'h1f, data_in[423:422],          {408{1'b0}},  8'h80};
                    667 : data_out = {data_in[1087:424],  5'h1f, data_in[423:421],          {408{1'b0}},  8'h80};
                    668 : data_out = {data_in[1087:424],  4'hf,  data_in[423:420],   8'h1,  {400{1'b0}},  8'h80};
                    669 : data_out = {data_in[1087:424],  3'h7,  data_in[423:419],   8'h3,  {400{1'b0}},  8'h80};
                    670 : data_out = {data_in[1087:424],  2'h3,  data_in[423:418],   8'h7,  {400{1'b0}},  8'h80};
                    671 : data_out = {data_in[1087:424],  1'h1,  data_in[423:417],   8'hf,  {400{1'b0}},  8'h80};
                    672 : data_out = {data_in[1087:416],                             8'h1f, {400{1'b0}},  8'h80};

                    673 : data_out = {data_in[1087:416],  7'h1f, data_in[415],              {400{1'b0}},  8'h80};
                    674 : data_out = {data_in[1087:416],  6'h1f, data_in[415:414],          {400{1'b0}},  8'h80};
                    675 : data_out = {data_in[1087:416],  5'h1f, data_in[415:413],          {400{1'b0}},  8'h80};
                    676 : data_out = {data_in[1087:416],  4'hf,  data_in[415:412],   8'h1,  {392{1'b0}},  8'h80};
                    677 : data_out = {data_in[1087:416],  3'h7,  data_in[415:411],   8'h3,  {392{1'b0}},  8'h80};
                    678 : data_out = {data_in[1087:416],  2'h3,  data_in[415:410],   8'h7,  {392{1'b0}},  8'h80};
                    679 : data_out = {data_in[1087:416],  1'h1,  data_in[415:409],   8'hf,  {392{1'b0}},  8'h80};
                    680 : data_out = {data_in[1087:408],                             8'h1f, {392{1'b0}},  8'h80};

                    681 : data_out = {data_in[1087:408],  7'h1f, data_in[407],              {392{1'b0}},  8'h80};
                    682 : data_out = {data_in[1087:408],  6'h1f, data_in[407:406],          {392{1'b0}},  8'h80};
                    683 : data_out = {data_in[1087:408],  5'h1f, data_in[407:405],          {392{1'b0}},  8'h80};
                    684 : data_out = {data_in[1087:408],  4'hf,  data_in[407:404],   8'h1,  {384{1'b0}},  8'h80};
                    685 : data_out = {data_in[1087:408],  3'h7,  data_in[407:403],   8'h3,  {384{1'b0}},  8'h80};
                    686 : data_out = {data_in[1087:408],  2'h3,  data_in[407:402],   8'h7,  {384{1'b0}},  8'h80};
                    687 : data_out = {data_in[1087:408],  1'h1,  data_in[407:401],   8'hf,  {384{1'b0}},  8'h80};
                    688 : data_out = {data_in[1087:400],                             8'h1f, {384{1'b0}},  8'h80};

                    689 : data_out = {data_in[1087:400],  7'h1f, data_in[399],              {384{1'b0}},  8'h80};
                    690 : data_out = {data_in[1087:400],  6'h1f, data_in[399:398],          {384{1'b0}},  8'h80};
                    691 : data_out = {data_in[1087:400],  5'h1f, data_in[399:397],          {384{1'b0}},  8'h80};
                    692 : data_out = {data_in[1087:400],  4'hf,  data_in[399:396],   8'h1,  {376{1'b0}},  8'h80};
                    693 : data_out = {data_in[1087:400],  3'h7,  data_in[399:395],   8'h3,  {376{1'b0}},  8'h80};
                    694 : data_out = {data_in[1087:400],  2'h3,  data_in[399:394],   8'h7,  {376{1'b0}},  8'h80};
                    695 : data_out = {data_in[1087:400],  1'h1,  data_in[399:393],   8'hf,  {376{1'b0}},  8'h80};
                    696 : data_out = {data_in[1087:392],                             8'h1f, {376{1'b0}},  8'h80};

                    697 : data_out = {data_in[1087:392],  7'h1f, data_in[391],              {376{1'b0}},  8'h80};
                    698 : data_out = {data_in[1087:392],  6'h1f, data_in[391:390],          {376{1'b0}},  8'h80};
                    699 : data_out = {data_in[1087:392],  5'h1f, data_in[391:389],          {376{1'b0}},  8'h80};
                    700 : data_out = {data_in[1087:392],  4'hf,  data_in[391:388],   8'h1,  {368{1'b0}},  8'h80};
                    701 : data_out = {data_in[1087:392],  3'h7,  data_in[391:387],   8'h3,  {368{1'b0}},  8'h80};
                    702 : data_out = {data_in[1087:392],  2'h3,  data_in[391:386],   8'h7,  {368{1'b0}},  8'h80};
                    703 : data_out = {data_in[1087:392],  1'h1,  data_in[391:385],   8'hf,  {368{1'b0}},  8'h80};
                    704 : data_out = {data_in[1087:384],                             8'h1f, {368{1'b0}},  8'h80};

                    705 : data_out = {data_in[1087:384],  7'h1f, data_in[383],              {368{1'b0}},  8'h80};
                    706 : data_out = {data_in[1087:384],  6'h1f, data_in[383:382],          {368{1'b0}},  8'h80};
                    707 : data_out = {data_in[1087:384],  5'h1f, data_in[383:381],          {368{1'b0}},  8'h80};
                    708 : data_out = {data_in[1087:384],  4'hf,  data_in[383:380],   8'h1,  {360{1'b0}},  8'h80};
                    709 : data_out = {data_in[1087:384],  3'h7,  data_in[383:379],   8'h3,  {360{1'b0}},  8'h80};
                    710 : data_out = {data_in[1087:384],  2'h3,  data_in[383:378],   8'h7,  {360{1'b0}},  8'h80};
                    711 : data_out = {data_in[1087:384],  1'h1,  data_in[383:377],   8'hf,  {360{1'b0}},  8'h80};
                    712 : data_out = {data_in[1087:376],                             8'h1f, {360{1'b0}},  8'h80};

                    713 : data_out = {data_in[1087:376],  7'h1f, data_in[375],              {360{1'b0}},  8'h80};
                    714 : data_out = {data_in[1087:376],  6'h1f, data_in[375:374],          {360{1'b0}},  8'h80};
                    715 : data_out = {data_in[1087:376],  5'h1f, data_in[375:373],          {360{1'b0}},  8'h80};
                    716 : data_out = {data_in[1087:376],  4'hf,  data_in[375:372],   8'h1,  {352{1'b0}},  8'h80};
                    717 : data_out = {data_in[1087:376],  3'h7,  data_in[375:371],   8'h3,  {352{1'b0}},  8'h80};
                    718 : data_out = {data_in[1087:376],  2'h3,  data_in[375:370],   8'h7,  {352{1'b0}},  8'h80};
                    719 : data_out = {data_in[1087:376],  1'h1,  data_in[375:369],   8'hf,  {352{1'b0}},  8'h80};
                    720 : data_out = {data_in[1087:368],                             8'h1f, {352{1'b0}},  8'h80};

                    721 : data_out = {data_in[1087:368],  7'h1f, data_in[367],              {352{1'b0}},  8'h80};
                    722 : data_out = {data_in[1087:368],  6'h1f, data_in[367:366],          {352{1'b0}},  8'h80};
                    723 : data_out = {data_in[1087:368],  5'h1f, data_in[367:365],          {352{1'b0}},  8'h80};
                    724 : data_out = {data_in[1087:368],  4'hf,  data_in[367:364],   8'h1,  {344{1'b0}},  8'h80};
                    725 : data_out = {data_in[1087:368],  3'h7,  data_in[367:363],   8'h3,  {344{1'b0}},  8'h80};
                    726 : data_out = {data_in[1087:368],  2'h3,  data_in[367:362],   8'h7,  {344{1'b0}},  8'h80};
                    727 : data_out = {data_in[1087:368],  1'h1,  data_in[367:361],   8'hf,  {344{1'b0}},  8'h80};
                    728 : data_out = {data_in[1087:360],                             8'h1f, {344{1'b0}},  8'h80};

                    729 : data_out = {data_in[1087:360],  7'h1f, data_in[359],              {344{1'b0}},  8'h80};
                    730 : data_out = {data_in[1087:360],  6'h1f, data_in[359:358],          {344{1'b0}},  8'h80};
                    731 : data_out = {data_in[1087:360],  5'h1f, data_in[359:357],          {344{1'b0}},  8'h80};
                    732 : data_out = {data_in[1087:360],  4'hf,  data_in[359:356],   8'h1,  {336{1'b0}},  8'h80};
                    733 : data_out = {data_in[1087:360],  3'h7,  data_in[359:355],   8'h3,  {336{1'b0}},  8'h80};
                    734 : data_out = {data_in[1087:360],  2'h3,  data_in[359:354],   8'h7,  {336{1'b0}},  8'h80};
                    735 : data_out = {data_in[1087:360],  1'h1,  data_in[359:353],   8'hf,  {336{1'b0}},  8'h80};
                    736 : data_out = {data_in[1087:352],                             8'h1f, {336{1'b0}},  8'h80};

                    737 : data_out = {data_in[1087:352],  7'h1f, data_in[351],              {336{1'b0}},  8'h80};
                    738 : data_out = {data_in[1087:352],  6'h1f, data_in[351:350],          {336{1'b0}},  8'h80};
                    739 : data_out = {data_in[1087:352],  5'h1f, data_in[351:349],          {336{1'b0}},  8'h80};
                    740 : data_out = {data_in[1087:352],  4'hf,  data_in[351:348],   8'h1,  {328{1'b0}},  8'h80};
                    741 : data_out = {data_in[1087:352],  3'h7,  data_in[351:347],   8'h3,  {328{1'b0}},  8'h80};
                    742 : data_out = {data_in[1087:352],  2'h3,  data_in[351:346],   8'h7,  {328{1'b0}},  8'h80};
                    743 : data_out = {data_in[1087:352],  1'h1,  data_in[351:345],   8'hf,  {328{1'b0}},  8'h80};
                    744 : data_out = {data_in[1087:344],                             8'h1f, {328{1'b0}},  8'h80};

                    745 : data_out = {data_in[1087:344],  7'h1f, data_in[343],              {328{1'b0}},  8'h80};
                    746 : data_out = {data_in[1087:344],  6'h1f, data_in[343:342],          {328{1'b0}},  8'h80};
                    747 : data_out = {data_in[1087:344],  5'h1f, data_in[343:341],          {328{1'b0}},  8'h80};
                    748 : data_out = {data_in[1087:344],  4'hf,  data_in[343:340],   8'h1,  {320{1'b0}},  8'h80};
                    749 : data_out = {data_in[1087:344],  3'h7,  data_in[343:339],   8'h3,  {320{1'b0}},  8'h80};
                    750 : data_out = {data_in[1087:344],  2'h3,  data_in[343:338],   8'h7,  {320{1'b0}},  8'h80};
                    751 : data_out = {data_in[1087:344],  1'h1,  data_in[343:337],   8'hf,  {320{1'b0}},  8'h80};
                    752 : data_out = {data_in[1087:336],                             8'h1f, {320{1'b0}},  8'h80};

                    753 : data_out = {data_in[1087:336],  7'h1f, data_in[335],              {320{1'b0}},  8'h80};
                    754 : data_out = {data_in[1087:336],  6'h1f, data_in[335:334],          {320{1'b0}},  8'h80};
                    755 : data_out = {data_in[1087:336],  5'h1f, data_in[335:333],          {320{1'b0}},  8'h80};
                    756 : data_out = {data_in[1087:336],  4'hf,  data_in[335:332],   8'h1,  {312{1'b0}},  8'h80};
                    757 : data_out = {data_in[1087:336],  3'h7,  data_in[335:331],   8'h3,  {312{1'b0}},  8'h80};
                    758 : data_out = {data_in[1087:336],  2'h3,  data_in[335:330],   8'h7,  {312{1'b0}},  8'h80};
                    759 : data_out = {data_in[1087:336],  1'h1,  data_in[335:329],   8'hf,  {312{1'b0}},  8'h80};
                    760 : data_out = {data_in[1087:328],                             8'h1f, {312{1'b0}},  8'h80};

                    761 : data_out = {data_in[1087:328],  7'h1f, data_in[327],              {312{1'b0}},  8'h80};
                    762 : data_out = {data_in[1087:328],  6'h1f, data_in[327:326],          {312{1'b0}},  8'h80};
                    763 : data_out = {data_in[1087:328],  5'h1f, data_in[327:325],          {312{1'b0}},  8'h80};
                    764 : data_out = {data_in[1087:328],  4'hf,  data_in[327:324],   8'h1,  {304{1'b0}},  8'h80};
                    765 : data_out = {data_in[1087:328],  3'h7,  data_in[327:323],   8'h3,  {304{1'b0}},  8'h80};
                    766 : data_out = {data_in[1087:328],  2'h3,  data_in[327:322],   8'h7,  {304{1'b0}},  8'h80};
                    767 : data_out = {data_in[1087:328],  1'h1,  data_in[327:321],   8'hf,  {304{1'b0}},  8'h80};
                    768 : data_out = {data_in[1087:320],                             8'h1f, {304{1'b0}},  8'h80};

                    769 : data_out = {data_in[1087:320],  7'h1f, data_in[319],              {304{1'b0}},  8'h80};
                    770 : data_out = {data_in[1087:320],  6'h1f, data_in[319:318],          {304{1'b0}},  8'h80};
                    771 : data_out = {data_in[1087:320],  5'h1f, data_in[319:317],          {304{1'b0}},  8'h80};
                    772 : data_out = {data_in[1087:320],  4'hf,  data_in[319:316],   8'h1,  {296{1'b0}},  8'h80};
                    773 : data_out = {data_in[1087:320],  3'h7,  data_in[319:315],   8'h3,  {296{1'b0}},  8'h80};
                    774 : data_out = {data_in[1087:320],  2'h3,  data_in[319:314],   8'h7,  {296{1'b0}},  8'h80};
                    775 : data_out = {data_in[1087:320],  1'h1,  data_in[319:313],   8'hf,  {296{1'b0}},  8'h80};
                    776 : data_out = {data_in[1087:312],                             8'h1f, {296{1'b0}},  8'h80};

                    777 : data_out = {data_in[1087:312],  7'h1f, data_in[311],              {296{1'b0}},  8'h80};
                    778 : data_out = {data_in[1087:312],  6'h1f, data_in[311:310],          {296{1'b0}},  8'h80};
                    779 : data_out = {data_in[1087:312],  5'h1f, data_in[311:309],          {296{1'b0}},  8'h80};
                    780 : data_out = {data_in[1087:312],  4'hf,  data_in[311:308],   8'h1,  {288{1'b0}},  8'h80};
                    781 : data_out = {data_in[1087:312],  3'h7,  data_in[311:307],   8'h3,  {288{1'b0}},  8'h80};
                    782 : data_out = {data_in[1087:312],  2'h3,  data_in[311:306],   8'h7,  {288{1'b0}},  8'h80};
                    783 : data_out = {data_in[1087:312],  1'h1,  data_in[311:305],   8'hf,  {288{1'b0}},  8'h80};
                    784 : data_out = {data_in[1087:304],                             8'h1f, {288{1'b0}},  8'h80};

                    785 : data_out = {data_in[1087:304],  7'h1f, data_in[303],              {288{1'b0}},  8'h80};
                    786 : data_out = {data_in[1087:304],  6'h1f, data_in[303:302],          {288{1'b0}},  8'h80};
                    787 : data_out = {data_in[1087:304],  5'h1f, data_in[303:301],          {288{1'b0}},  8'h80};
                    788 : data_out = {data_in[1087:304],  4'hf,  data_in[303:300],   8'h1,  {280{1'b0}},  8'h80};
                    789 : data_out = {data_in[1087:304],  3'h7,  data_in[303:299],   8'h3,  {280{1'b0}},  8'h80};
                    790 : data_out = {data_in[1087:304],  2'h3,  data_in[303:298],   8'h7,  {280{1'b0}},  8'h80};
                    791 : data_out = {data_in[1087:304],  1'h1,  data_in[303:297],   8'hf,  {280{1'b0}},  8'h80};
                    792 : data_out = {data_in[1087:296],                             8'h1f, {280{1'b0}},  8'h80};

                    793 : data_out = {data_in[1087:296],  7'h1f, data_in[295],              {280{1'b0}},  8'h80};
                    794 : data_out = {data_in[1087:296],  6'h1f, data_in[295:294],          {280{1'b0}},  8'h80};
                    795 : data_out = {data_in[1087:296],  5'h1f, data_in[295:293],          {280{1'b0}},  8'h80};
                    796 : data_out = {data_in[1087:296],  4'hf,  data_in[295:292],   8'h1,  {272{1'b0}},  8'h80};
                    797 : data_out = {data_in[1087:296],  3'h7,  data_in[295:291],   8'h3,  {272{1'b0}},  8'h80};
                    798 : data_out = {data_in[1087:296],  2'h3,  data_in[295:290],   8'h7,  {272{1'b0}},  8'h80};
                    799 : data_out = {data_in[1087:296],  1'h1,  data_in[295:289],   8'hf,  {272{1'b0}},  8'h80};
                    800 : data_out = {data_in[1087:288],                             8'h1f, {272{1'b0}},  8'h80};

                    801 : data_out = {data_in[1087:288],  7'h1f, data_in[287],              {272{1'b0}},  8'h80};
                    802 : data_out = {data_in[1087:288],  6'h1f, data_in[287:286],          {272{1'b0}},  8'h80};
                    803 : data_out = {data_in[1087:288],  5'h1f, data_in[287:285],          {272{1'b0}},  8'h80};
                    804 : data_out = {data_in[1087:288],  4'hf,  data_in[287:284],   8'h1,  {264{1'b0}},  8'h80};
                    805 : data_out = {data_in[1087:288],  3'h7,  data_in[287:283],   8'h3,  {264{1'b0}},  8'h80};
                    806 : data_out = {data_in[1087:288],  2'h3,  data_in[287:282],   8'h7,  {264{1'b0}},  8'h80};
                    807 : data_out = {data_in[1087:288],  1'h1,  data_in[287:281],   8'hf,  {264{1'b0}},  8'h80};
                    808 : data_out = {data_in[1087:280],                             8'h1f, {264{1'b0}},  8'h80};

                    809 : data_out = {data_in[1087:280],  7'h1f, data_in[279],              {264{1'b0}},  8'h80};
                    810 : data_out = {data_in[1087:280],  6'h1f, data_in[279:278],          {264{1'b0}},  8'h80};
                    811 : data_out = {data_in[1087:280],  5'h1f, data_in[279:277],          {264{1'b0}},  8'h80};
                    812 : data_out = {data_in[1087:280],  4'hf,  data_in[279:276],   8'h1,  {256{1'b0}},  8'h80};
                    813 : data_out = {data_in[1087:280],  3'h7,  data_in[279:275],   8'h3,  {256{1'b0}},  8'h80};
                    814 : data_out = {data_in[1087:280],  2'h3,  data_in[279:274],   8'h7,  {256{1'b0}},  8'h80};
                    815 : data_out = {data_in[1087:280],  1'h1,  data_in[279:273],   8'hf,  {256{1'b0}},  8'h80};
                    816 : data_out = {data_in[1087:272],                             8'h1f, {256{1'b0}},  8'h80};

                    817 : data_out = {data_in[1087:272],  7'h1f, data_in[271],              {256{1'b0}},  8'h80};
                    818 : data_out = {data_in[1087:272],  6'h1f, data_in[271:270],          {256{1'b0}},  8'h80};
                    819 : data_out = {data_in[1087:272],  5'h1f, data_in[271:269],          {256{1'b0}},  8'h80};
                    820 : data_out = {data_in[1087:272],  4'hf,  data_in[271:268],   8'h1,  {248{1'b0}},  8'h80};
                    821 : data_out = {data_in[1087:272],  3'h7,  data_in[271:267],   8'h3,  {248{1'b0}},  8'h80};
                    822 : data_out = {data_in[1087:272],  2'h3,  data_in[271:266],   8'h7,  {248{1'b0}},  8'h80};
                    823 : data_out = {data_in[1087:272],  1'h1,  data_in[271:265],   8'hf,  {248{1'b0}},  8'h80};
                    824 : data_out = {data_in[1087:264],                             8'h1f, {248{1'b0}},  8'h80};

                    825 : data_out = {data_in[1087:264],  7'h1f, data_in[263],              {248{1'b0}},  8'h80};
                    826 : data_out = {data_in[1087:264],  6'h1f, data_in[263:262],          {248{1'b0}},  8'h80};
                    827 : data_out = {data_in[1087:264],  5'h1f, data_in[263:261],          {248{1'b0}},  8'h80};
                    828 : data_out = {data_in[1087:264],  4'hf,  data_in[263:260],   8'h1,  {240{1'b0}},  8'h80};
                    829 : data_out = {data_in[1087:264],  3'h7,  data_in[263:259],   8'h3,  {240{1'b0}},  8'h80};
                    830 : data_out = {data_in[1087:264],  2'h3,  data_in[263:258],   8'h7,  {240{1'b0}},  8'h80};
                    831 : data_out = {data_in[1087:264],  1'h1,  data_in[263:257],   8'hf,  {240{1'b0}},  8'h80};
                    832 : data_out = {data_in[1087:256],                             8'h1f, {240{1'b0}},  8'h80};

                    833 : data_out = {data_in[1087:256],  7'h1f, data_in[255],              {240{1'b0}},  8'h80};
                    834 : data_out = {data_in[1087:256],  6'h1f, data_in[255:254],          {240{1'b0}},  8'h80};
                    835 : data_out = {data_in[1087:256],  5'h1f, data_in[255:253],          {240{1'b0}},  8'h80};
                    836 : data_out = {data_in[1087:256],  4'hf,  data_in[255:252],   8'h1,  {232{1'b0}},  8'h80};
                    837 : data_out = {data_in[1087:256],  3'h7,  data_in[255:251],   8'h3,  {232{1'b0}},  8'h80};
                    838 : data_out = {data_in[1087:256],  2'h3,  data_in[255:250],   8'h7,  {232{1'b0}},  8'h80};
                    839 : data_out = {data_in[1087:256],  1'h1,  data_in[255:249],   8'hf,  {232{1'b0}},  8'h80};
                    840 : data_out = {data_in[1087:248],                             8'h1f, {232{1'b0}},  8'h80};

                    841 : data_out = {data_in[1087:248],  7'h1f, data_in[247],              {232{1'b0}},  8'h80};
                    842 : data_out = {data_in[1087:248],  6'h1f, data_in[247:246],          {232{1'b0}},  8'h80};
                    843 : data_out = {data_in[1087:248],  5'h1f, data_in[247:245],          {232{1'b0}},  8'h80};
                    844 : data_out = {data_in[1087:248],  4'hf,  data_in[247:244],   8'h1,  {224{1'b0}},  8'h80};
                    845 : data_out = {data_in[1087:248],  3'h7,  data_in[247:243],   8'h3,  {224{1'b0}},  8'h80};
                    846 : data_out = {data_in[1087:248],  2'h3,  data_in[247:242],   8'h7,  {224{1'b0}},  8'h80};
                    847 : data_out = {data_in[1087:248],  1'h1,  data_in[247:241],   8'hf,  {224{1'b0}},  8'h80};
                    848 : data_out = {data_in[1087:240],                             8'h1f, {224{1'b0}},  8'h80};

                    849 : data_out = {data_in[1087:240],  7'h1f, data_in[239],              {224{1'b0}},  8'h80};
                    850 : data_out = {data_in[1087:240],  6'h1f, data_in[239:238],          {224{1'b0}},  8'h80};
                    851 : data_out = {data_in[1087:240],  5'h1f, data_in[239:237],          {224{1'b0}},  8'h80};
                    852 : data_out = {data_in[1087:240],  4'hf,  data_in[239:236],   8'h1,  {216{1'b0}},  8'h80};
                    853 : data_out = {data_in[1087:240],  3'h7,  data_in[239:235],   8'h3,  {216{1'b0}},  8'h80};
                    854 : data_out = {data_in[1087:240],  2'h3,  data_in[239:234],   8'h7,  {216{1'b0}},  8'h80};
                    855 : data_out = {data_in[1087:240],  1'h1,  data_in[239:233],   8'hf,  {216{1'b0}},  8'h80};
                    856 : data_out = {data_in[1087:232],                             8'h1f, {216{1'b0}},  8'h80};

                    857 : data_out = {data_in[1087:232],  7'h1f, data_in[231],              {216{1'b0}},  8'h80};
                    858 : data_out = {data_in[1087:232],  6'h1f, data_in[231:230],          {216{1'b0}},  8'h80};
                    859 : data_out = {data_in[1087:232],  5'h1f, data_in[231:229],          {216{1'b0}},  8'h80};
                    860 : data_out = {data_in[1087:232],  4'hf,  data_in[231:228],   8'h1,  {208{1'b0}},  8'h80};
                    861 : data_out = {data_in[1087:232],  3'h7,  data_in[231:227],   8'h3,  {208{1'b0}},  8'h80};
                    862 : data_out = {data_in[1087:232],  2'h3,  data_in[231:226],   8'h7,  {208{1'b0}},  8'h80};
                    863 : data_out = {data_in[1087:232],  1'h1,  data_in[231:225],   8'hf,  {208{1'b0}},  8'h80};
                    864 : data_out = {data_in[1087:224],                             8'h1f, {208{1'b0}},  8'h80};

                    865 : data_out = {data_in[1087:224],  7'h1f, data_in[223],              {208{1'b0}},  8'h80};
                    866 : data_out = {data_in[1087:224],  6'h1f, data_in[223:222],          {208{1'b0}},  8'h80};
                    867 : data_out = {data_in[1087:224],  5'h1f, data_in[223:221],          {208{1'b0}},  8'h80};
                    868 : data_out = {data_in[1087:224],  4'hf,  data_in[223:220],   8'h1,  {200{1'b0}},  8'h80};
                    869 : data_out = {data_in[1087:224],  3'h7,  data_in[223:219],   8'h3,  {200{1'b0}},  8'h80};
                    870 : data_out = {data_in[1087:224],  2'h3,  data_in[223:218],   8'h7,  {200{1'b0}},  8'h80};
                    871 : data_out = {data_in[1087:224],  1'h1,  data_in[223:217],   8'hf,  {200{1'b0}},  8'h80};
                    872 : data_out = {data_in[1087:216],                             8'h1f, {200{1'b0}},  8'h80};

                    873 : data_out = {data_in[1087:216],  7'h1f, data_in[215],              {200{1'b0}},  8'h80};
                    874 : data_out = {data_in[1087:216],  6'h1f, data_in[215:214],          {200{1'b0}},  8'h80};
                    875 : data_out = {data_in[1087:216],  5'h1f, data_in[215:213],          {200{1'b0}},  8'h80};
                    876 : data_out = {data_in[1087:216],  4'hf,  data_in[215:212],   8'h1,  {192{1'b0}},  8'h80};
                    877 : data_out = {data_in[1087:216],  3'h7,  data_in[215:211],   8'h3,  {192{1'b0}},  8'h80};
                    878 : data_out = {data_in[1087:216],  2'h3,  data_in[215:210],   8'h7,  {192{1'b0}},  8'h80};
                    879 : data_out = {data_in[1087:216],  1'h1,  data_in[215:209],   8'hf,  {192{1'b0}},  8'h80};
                    880 : data_out = {data_in[1087:208],                             8'h1f, {192{1'b0}},  8'h80};

                    881 : data_out = {data_in[1087:208],  7'h1f, data_in[207],              {192{1'b0}},  8'h80};
                    882 : data_out = {data_in[1087:208],  6'h1f, data_in[207:206],          {192{1'b0}},  8'h80};
                    883 : data_out = {data_in[1087:208],  5'h1f, data_in[207:205],          {192{1'b0}},  8'h80};
                    884 : data_out = {data_in[1087:208],  4'hf,  data_in[207:204],   8'h1,  {184{1'b0}},  8'h80};
                    885 : data_out = {data_in[1087:208],  3'h7,  data_in[207:203],   8'h3,  {184{1'b0}},  8'h80};
                    886 : data_out = {data_in[1087:208],  2'h3,  data_in[207:202],   8'h7,  {184{1'b0}},  8'h80};
                    887 : data_out = {data_in[1087:208],  1'h1,  data_in[207:201],   8'hf,  {184{1'b0}},  8'h80};
                    888 : data_out = {data_in[1087:200],                             8'h1f, {184{1'b0}},  8'h80};

                    889 : data_out = {data_in[1087:200],  7'h1f, data_in[199],              {184{1'b0}},  8'h80};
                    890 : data_out = {data_in[1087:200],  6'h1f, data_in[199:198],          {184{1'b0}},  8'h80};
                    891 : data_out = {data_in[1087:200],  5'h1f, data_in[199:197],          {184{1'b0}},  8'h80};
                    892 : data_out = {data_in[1087:200],  4'hf,  data_in[199:196],   8'h1,  {176{1'b0}},  8'h80};
                    893 : data_out = {data_in[1087:200],  3'h7,  data_in[199:195],   8'h3,  {176{1'b0}},  8'h80};
                    894 : data_out = {data_in[1087:200],  2'h3,  data_in[199:194],   8'h7,  {176{1'b0}},  8'h80};
                    895 : data_out = {data_in[1087:200],  1'h1,  data_in[199:193],   8'hf,  {176{1'b0}},  8'h80};
                    896 : data_out = {data_in[1087:192],                             8'h1f, {176{1'b0}},  8'h80};

                    897 : data_out = {data_in[1087:192],  7'h1f, data_in[191],              {176{1'b0}},  8'h80};
                    898 : data_out = {data_in[1087:192],  6'h1f, data_in[191:190],          {176{1'b0}},  8'h80};
                    899 : data_out = {data_in[1087:192],  5'h1f, data_in[191:189],          {176{1'b0}},  8'h80};
                    900 : data_out = {data_in[1087:192],  4'hf,  data_in[191:188],   8'h1,  {168{1'b0}},  8'h80};
                    901 : data_out = {data_in[1087:192],  3'h7,  data_in[191:187],   8'h3,  {168{1'b0}},  8'h80};
                    902 : data_out = {data_in[1087:192],  2'h3,  data_in[191:186],   8'h7,  {168{1'b0}},  8'h80};
                    903 : data_out = {data_in[1087:192],  1'h1,  data_in[191:185],   8'hf,  {168{1'b0}},  8'h80};
                    904 : data_out = {data_in[1087:184],                             8'h1f, {168{1'b0}},  8'h80};

                    905 : data_out = {data_in[1087:184],  7'h1f, data_in[183],              {168{1'b0}},  8'h80};
                    906 : data_out = {data_in[1087:184],  6'h1f, data_in[183:182],          {168{1'b0}},  8'h80};
                    907 : data_out = {data_in[1087:184],  5'h1f, data_in[183:181],          {168{1'b0}},  8'h80};
                    908 : data_out = {data_in[1087:184],  4'hf,  data_in[183:180],   8'h1,  {160{1'b0}},  8'h80};
                    909 : data_out = {data_in[1087:184],  3'h7,  data_in[183:179],   8'h3,  {160{1'b0}},  8'h80};
                    910 : data_out = {data_in[1087:184],  2'h3,  data_in[183:178],   8'h7,  {160{1'b0}},  8'h80};
                    911 : data_out = {data_in[1087:184],  1'h1,  data_in[183:177],   8'hf,  {160{1'b0}},  8'h80};
                    912 : data_out = {data_in[1087:176],                             8'h1f, {160{1'b0}},  8'h80};

                    913 : data_out = {data_in[1087:176],  7'h1f, data_in[175],              {160{1'b0}},  8'h80};
                    914 : data_out = {data_in[1087:176],  6'h1f, data_in[175:174],          {160{1'b0}},  8'h80};
                    915 : data_out = {data_in[1087:176],  5'h1f, data_in[175:173],          {160{1'b0}},  8'h80};
                    916 : data_out = {data_in[1087:176],  4'hf,  data_in[175:172],   8'h1,  {152{1'b0}},  8'h80};
                    917 : data_out = {data_in[1087:176],  3'h7,  data_in[175:171],   8'h3,  {152{1'b0}},  8'h80};
                    918 : data_out = {data_in[1087:176],  2'h3,  data_in[175:170],   8'h7,  {152{1'b0}},  8'h80};
                    919 : data_out = {data_in[1087:176],  1'h1,  data_in[175:169],   8'hf,  {152{1'b0}},  8'h80};
                    920 : data_out = {data_in[1087:168],                             8'h1f, {152{1'b0}},  8'h80};

                    921 : data_out = {data_in[1087:168],  7'h1f, data_in[167],              {152{1'b0}},  8'h80};
                    922 : data_out = {data_in[1087:168],  6'h1f, data_in[167:166],          {152{1'b0}},  8'h80};
                    923 : data_out = {data_in[1087:168],  5'h1f, data_in[167:165],          {152{1'b0}},  8'h80};
                    924 : data_out = {data_in[1087:168],  4'hf,  data_in[167:164],   8'h1,  {144{1'b0}},  8'h80};
                    925 : data_out = {data_in[1087:168],  3'h7,  data_in[167:163],   8'h3,  {144{1'b0}},  8'h80};
                    926 : data_out = {data_in[1087:168],  2'h3,  data_in[167:162],   8'h7,  {144{1'b0}},  8'h80};
                    927 : data_out = {data_in[1087:168],  1'h1,  data_in[167:161],   8'hf,  {144{1'b0}},  8'h80};
                    928 : data_out = {data_in[1087:160],                             8'h1f, {144{1'b0}},  8'h80};

                    929 : data_out = {data_in[1087:160],  7'h1f, data_in[159],              {144{1'b0}},  8'h80};
                    930 : data_out = {data_in[1087:160],  6'h1f, data_in[159:158],          {144{1'b0}},  8'h80};
                    931 : data_out = {data_in[1087:160],  5'h1f, data_in[159:157],          {144{1'b0}},  8'h80};
                    932 : data_out = {data_in[1087:160],  4'hf,  data_in[159:156],   8'h1,  {136{1'b0}},  8'h80};
                    933 : data_out = {data_in[1087:160],  3'h7,  data_in[159:155],   8'h3,  {136{1'b0}},  8'h80};
                    934 : data_out = {data_in[1087:160],  2'h3,  data_in[159:154],   8'h7,  {136{1'b0}},  8'h80};
                    935 : data_out = {data_in[1087:160],  1'h1,  data_in[159:153],   8'hf,  {136{1'b0}},  8'h80};
                    936 : data_out = {data_in[1087:152],                             8'h1f, {136{1'b0}},  8'h80};

                    937 : data_out = {data_in[1087:152],  7'h1f, data_in[151],              {136{1'b0}},  8'h80};
                    938 : data_out = {data_in[1087:152],  6'h1f, data_in[151:150],          {136{1'b0}},  8'h80};
                    939 : data_out = {data_in[1087:152],  5'h1f, data_in[151:149],          {136{1'b0}},  8'h80};
                    940 : data_out = {data_in[1087:152],  4'hf,  data_in[151:148],   8'h1,  {128{1'b0}},  8'h80};
                    941 : data_out = {data_in[1087:152],  3'h7,  data_in[151:147],   8'h3,  {128{1'b0}},  8'h80};
                    942 : data_out = {data_in[1087:152],  2'h3,  data_in[151:146],   8'h7,  {128{1'b0}},  8'h80};
                    943 : data_out = {data_in[1087:152],  1'h1,  data_in[151:145],   8'hf,  {128{1'b0}},  8'h80};
                    944 : data_out = {data_in[1087:144],                             8'h1f, {128{1'b0}},  8'h80};

                    945 : data_out = {data_in[1087:144],  7'h1f, data_in[143],              {128{1'b0}},  8'h80};
                    946 : data_out = {data_in[1087:144],  6'h1f, data_in[143:142],          {128{1'b0}},  8'h80};
                    947 : data_out = {data_in[1087:144],  5'h1f, data_in[143:141],          {128{1'b0}},  8'h80};
                    948 : data_out = {data_in[1087:144],  4'hf,  data_in[143:140],   8'h1,  {120{1'b0}},  8'h80};
                    949 : data_out = {data_in[1087:144],  3'h7,  data_in[143:139],   8'h3,  {120{1'b0}},  8'h80};
                    950 : data_out = {data_in[1087:144],  2'h3,  data_in[143:138],   8'h7,  {120{1'b0}},  8'h80};
                    951 : data_out = {data_in[1087:144],  1'h1,  data_in[143:137],   8'hf,  {120{1'b0}},  8'h80};
                    952 : data_out = {data_in[1087:136],                             8'h1f, {120{1'b0}},  8'h80};

                    953 : data_out = {data_in[1087:136],  7'h1f, data_in[135],              {120{1'b0}},  8'h80};
                    954 : data_out = {data_in[1087:136],  6'h1f, data_in[135:134],          {120{1'b0}},  8'h80};
                    955 : data_out = {data_in[1087:136],  5'h1f, data_in[135:133],          {120{1'b0}},  8'h80};
                    956 : data_out = {data_in[1087:136],  4'hf,  data_in[135:132],   8'h1,  {112{1'b0}},  8'h80};
                    957 : data_out = {data_in[1087:136],  3'h7,  data_in[135:131],   8'h3,  {112{1'b0}},  8'h80};
                    958 : data_out = {data_in[1087:136],  2'h3,  data_in[135:130],   8'h7,  {112{1'b0}},  8'h80};
                    959 : data_out = {data_in[1087:136],  1'h1,  data_in[135:129],   8'hf,  {112{1'b0}},  8'h80};
                    960 : data_out = {data_in[1087:128],                             8'h1f, {112{1'b0}},  8'h80};

                    961 : data_out = {data_in[1087:128],  7'h1f, data_in[127],              {112{1'b0}},  8'h80};
                    962 : data_out = {data_in[1087:128],  6'h1f, data_in[127:126],          {112{1'b0}},  8'h80};
                    963 : data_out = {data_in[1087:128],  5'h1f, data_in[127:125],          {112{1'b0}},  8'h80};
                    964 : data_out = {data_in[1087:128],  4'hf,  data_in[127:124],   8'h1,  {104{1'b0}},  8'h80};
                    965 : data_out = {data_in[1087:128],  3'h7,  data_in[127:123],   8'h3,  {104{1'b0}},  8'h80};
                    966 : data_out = {data_in[1087:128],  2'h3,  data_in[127:122],   8'h7,  {104{1'b0}},  8'h80};
                    967 : data_out = {data_in[1087:128],  1'h1,  data_in[127:121],   8'hf,  {104{1'b0}},  8'h80};
                    968 : data_out = {data_in[1087:120],                             8'h1f, {104{1'b0}},  8'h80};

                    969 : data_out = {data_in[1087:120],  7'h1f, data_in[119],              {104{1'b0}},  8'h80};
                    970 : data_out = {data_in[1087:120],  6'h1f, data_in[119:118],          {104{1'b0}},  8'h80};
                    971 : data_out = {data_in[1087:120],  5'h1f, data_in[119:117],          {104{1'b0}},  8'h80};
                    972 : data_out = {data_in[1087:120],  4'hf,  data_in[119:116],   8'h1,  {96{1'b0}},   8'h80};
                    973 : data_out = {data_in[1087:120],  3'h7,  data_in[119:115],   8'h3,  {96{1'b0}},   8'h80};
                    974 : data_out = {data_in[1087:120],  2'h3,  data_in[119:114],   8'h7,  {96{1'b0}},   8'h80};
                    975 : data_out = {data_in[1087:120],  1'h1,  data_in[119:113],   8'hf,  {96{1'b0}},   8'h80};
                    976 : data_out = {data_in[1087:112],                             8'h1f, {96{1'b0}},   8'h80};

                    977 : data_out = {data_in[1087:112],  7'h1f, data_in[111],              {96{1'b0}},   8'h80};
                    978 : data_out = {data_in[1087:112],  6'h1f, data_in[111:110],          {96{1'b0}},   8'h80};
                    979 : data_out = {data_in[1087:112],  5'h1f, data_in[111:109],          {96{1'b0}},   8'h80};
                    980 : data_out = {data_in[1087:112],  4'hf,  data_in[111:108],   8'h1,  {88{1'b0}},   8'h80};
                    981 : data_out = {data_in[1087:112],  3'h7,  data_in[111:107],   8'h3,  {88{1'b0}},   8'h80};
                    982 : data_out = {data_in[1087:112],  2'h3,  data_in[111:106],   8'h7,  {88{1'b0}},   8'h80};
                    983 : data_out = {data_in[1087:112],  1'h1,  data_in[111:105],   8'hf,  {88{1'b0}},   8'h80};
                    984 : data_out = {data_in[1087:104],                             8'h1f, {88{1'b0}},   8'h80};

                    985 : data_out = {data_in[1087:104],  7'h1f, data_in[103],              {88{1'b0}},   8'h80};
                    986 : data_out = {data_in[1087:104],  6'h1f, data_in[103:102],          {88{1'b0}},   8'h80};
                    987 : data_out = {data_in[1087:104],  5'h1f, data_in[103:101],          {88{1'b0}},   8'h80};
                    988 : data_out = {data_in[1087:104],  4'hf,  data_in[103:100],   8'h1,  {80{1'b0}},   8'h80};
                    989 : data_out = {data_in[1087:104],  3'h7,  data_in[103:99],    8'h3,  {80{1'b0}},   8'h80};
                    990 : data_out = {data_in[1087:104],  2'h3,  data_in[103:98],    8'h7,  {80{1'b0}},   8'h80};
                    991 : data_out = {data_in[1087:104],  1'h1,  data_in[103:97],    8'hf,  {80{1'b0}},   8'h80};
                    992 : data_out = {data_in[1087:96],                              8'h1f, {80{1'b0}},   8'h80};

                    993 : data_out = {data_in[1087:96],   7'h1f, data_in[95],               {80{1'b0}},   8'h80};
                    994 : data_out = {data_in[1087:96],   6'h1f, data_in[95:94],            {80{1'b0}},   8'h80};
                    995 : data_out = {data_in[1087:96],   5'h1f, data_in[95:93],            {80{1'b0}},   8'h80};
                    996 : data_out = {data_in[1087:96],   4'hf,  data_in[95:92],     8'h1,  {72{1'b0}},   8'h80};
                    997 : data_out = {data_in[1087:96],   3'h7,  data_in[95:91],     8'h3,  {72{1'b0}},   8'h80};
                    998 : data_out = {data_in[1087:96],   2'h3,  data_in[95:90],     8'h7,  {72{1'b0}},   8'h80};
                    999 : data_out = {data_in[1087:96],   1'h1,  data_in[95:89],     8'hf,  {72{1'b0}},   8'h80};
                    1000: data_out = {data_in[1087:88],                              8'h1f, {72{1'b0}},   8'h80};

                    1001: data_out = {data_in[1087:88],   7'h1f, data_in[87],               {72{1'b0}},   8'h80};
                    1002: data_out = {data_in[1087:88],   6'h1f, data_in[87:86],            {72{1'b0}},   8'h80};
                    1003: data_out = {data_in[1087:88],   5'h1f, data_in[87:85],            {72{1'b0}},   8'h80};
                    1004: data_out = {data_in[1087:88],   4'hf,  data_in[87:84],     8'h1,  {64{1'b0}},   8'h80};
                    1005: data_out = {data_in[1087:88],   3'h7,  data_in[87:83],     8'h3,  {64{1'b0}},   8'h80};
                    1006: data_out = {data_in[1087:88],   2'h3,  data_in[87:82],     8'h7,  {64{1'b0}},   8'h80};
                    1007: data_out = {data_in[1087:88],   1'h1,  data_in[87:81],     8'hf,  {64{1'b0}},   8'h80};
                    1008: data_out = {data_in[1087:80],                              8'h1f, {64{1'b0}},   8'h80};

                    1009: data_out = {data_in[1087:80],   7'h1f, data_in[79],               {64{1'b0}},   8'h80};
                    1010: data_out = {data_in[1087:80],   6'h1f, data_in[79:78],            {64{1'b0}},   8'h80};
                    1011: data_out = {data_in[1087:80],   5'h1f, data_in[79:77],            {64{1'b0}},   8'h80};
                    1012: data_out = {data_in[1087:80],   4'hf,  data_in[79:76],     8'h1,  {56{1'b0}},   8'h80};
                    1013: data_out = {data_in[1087:80],   3'h7,  data_in[79:75],     8'h3,  {56{1'b0}},   8'h80};
                    1014: data_out = {data_in[1087:80],   2'h3,  data_in[79:74],     8'h7,  {56{1'b0}},   8'h80};
                    1015: data_out = {data_in[1087:80],   1'h1,  data_in[79:73],     8'hf,  {56{1'b0}},   8'h80};
                    1016: data_out = {data_in[1087:72],                              8'h1f, {56{1'b0}},   8'h80};

                    1017: data_out = {data_in[1087:72],   7'h1f, data_in[71],               {56{1'b0}},   8'h80};
                    1018: data_out = {data_in[1087:72],   6'h1f, data_in[71:70],            {56{1'b0}},   8'h80};
                    1019: data_out = {data_in[1087:72],   5'h1f, data_in[71:69],            {56{1'b0}},   8'h80};
                    1020: data_out = {data_in[1087:72],   4'hf,  data_in[71:68],     8'h1,  {48{1'b0}},   8'h80};
                    1021: data_out = {data_in[1087:72],   3'h7,  data_in[71:67],     8'h3,  {48{1'b0}},   8'h80};
                    1022: data_out = {data_in[1087:72],   2'h3,  data_in[71:66],     8'h7,  {48{1'b0}},   8'h80};
                    1023: data_out = {data_in[1087:72],   1'h1,  data_in[71:65],     8'hf,  {48{1'b0}},   8'h80};
                    1024: data_out = {data_in[1087:64],                              8'h1f, {48{1'b0}},   8'h80};

                    1025: data_out = {data_in[1087:64],   7'h1f, data_in[63],               {48{1'b0}},   8'h80};
                    1026: data_out = {data_in[1087:64],   6'h1f, data_in[63:62],            {48{1'b0}},   8'h80};
                    1027: data_out = {data_in[1087:64],   5'h1f, data_in[63:61],            {48{1'b0}},   8'h80};
                    1028: data_out = {data_in[1087:64],   4'hf,  data_in[63:60],     8'h1,  {40{1'b0}},   8'h80};
                    1029: data_out = {data_in[1087:64],   3'h7,  data_in[63:59],     8'h3,  {40{1'b0}},   8'h80};
                    1030: data_out = {data_in[1087:64],   2'h3,  data_in[63:58],     8'h7,  {40{1'b0}},   8'h80};
                    1031: data_out = {data_in[1087:64],   1'h1,  data_in[63:57],     8'hf,  {40{1'b0}},   8'h80};
                    1032: data_out = {data_in[1087:56],                              8'h1f, {40{1'b0}},   8'h80};

                    1033: data_out = {data_in[1087:56],   7'h1f, data_in[55],               {40{1'b0}},   8'h80};
                    1034: data_out = {data_in[1087:56],   6'h1f, data_in[55:54],            {40{1'b0}},   8'h80};
                    1035: data_out = {data_in[1087:56],   5'h1f, data_in[55:53],            {40{1'b0}},   8'h80};
                    1036: data_out = {data_in[1087:56],   4'hf,  data_in[55:52],     8'h1,  {32{1'b0}},   8'h80};
                    1037: data_out = {data_in[1087:56],   3'h7,  data_in[55:51],     8'h3,  {32{1'b0}},   8'h80};
                    1038: data_out = {data_in[1087:56],   2'h3,  data_in[55:50],     8'h7,  {32{1'b0}},   8'h80};
                    1039: data_out = {data_in[1087:56],   1'h1,  data_in[55:49],     8'hf,  {32{1'b0}},   8'h80};
                    1040: data_out = {data_in[1087:48],                              8'h1f, {32{1'b0}},   8'h80};

                    1041: data_out = {data_in[1087:48],   7'h1f, data_in[47],               {32{1'b0}},   8'h80};
                    1042: data_out = {data_in[1087:48],   6'h1f, data_in[47:46],            {32{1'b0}},   8'h80};
                    1043: data_out = {data_in[1087:48],   5'h1f, data_in[47:45],            {32{1'b0}},   8'h80};
                    1044: data_out = {data_in[1087:48],   4'hf,  data_in[47:44],     8'h1,  {24{1'b0}},   8'h80};
                    1045: data_out = {data_in[1087:48],   3'h7,  data_in[47:43],     8'h3,  {24{1'b0}},   8'h80};
                    1046: data_out = {data_in[1087:48],   2'h3,  data_in[47:42],     8'h7,  {24{1'b0}},   8'h80};
                    1047: data_out = {data_in[1087:48],   1'h1,  data_in[47:41],     8'hf,  {24{1'b0}},   8'h80};
                    1048: data_out = {data_in[1087:40],                              8'h1f, {24{1'b0}},   8'h80};

                    1049: data_out = {data_in[1087:40],   7'h1f, data_in[39],               {24{1'b0}},   8'h80};
                    1050: data_out = {data_in[1087:40],   6'h1f, data_in[39:38],            {24{1'b0}},   8'h80};
                    1051: data_out = {data_in[1087:40],   5'h1f, data_in[39:37],            {24{1'b0}},   8'h80};
                    1052: data_out = {data_in[1087:40],   4'hf,  data_in[39:36],     8'h1,  {16{1'b0}},   8'h80};
                    1053: data_out = {data_in[1087:40],   3'h7,  data_in[39:35],     8'h3,  {16{1'b0}},   8'h80};
                    1054: data_out = {data_in[1087:40],   2'h3,  data_in[39:34],     8'h7,  {16{1'b0}},   8'h80};
                    1055: data_out = {data_in[1087:40],   1'h1,  data_in[39:33],     8'hf,  {16{1'b0}},   8'h80};
                    1056: data_out = {data_in[1087:32],                              8'h1f, {16{1'b0}},   8'h80};

                    1057: data_out = {data_in[1087:32],   7'h1f, data_in[31],               {16{1'b0}},   8'h80};
                    1058: data_out = {data_in[1087:32],   6'h1f, data_in[31:30],            {16{1'b0}},   8'h80};
                    1059: data_out = {data_in[1087:32],   5'h1f, data_in[31:29],            {16{1'b0}},   8'h80};
                    1060: data_out = {data_in[1087:32],   4'hf,  data_in[31:28],     8'h1,  {8{1'b0}},    8'h80};
                    1061: data_out = {data_in[1087:32],   3'h7,  data_in[31:27],     8'h3,  {8{1'b0}},    8'h80};
                    1062: data_out = {data_in[1087:32],   2'h3,  data_in[31:26],     8'h7,  {8{1'b0}},    8'h80};
                    1063: data_out = {data_in[1087:32],   1'h1,  data_in[31:25],     8'hf,  {8{1'b0}},    8'h80};
                    1064: data_out = {data_in[1087:24],                              8'h1f, {8{1'b0}},    8'h80};

                    1065: data_out = {data_in[1087:24],   7'h1f, data_in[23],               {8{1'b0}},    8'h80};
                    1066: data_out = {data_in[1087:24],   6'h1f, data_in[23:22],            {8{1'b0}},    8'h80};
                    1067: data_out = {data_in[1087:24],   5'h1f, data_in[23:21],            {8{1'b0}},    8'h80};
                    1068: data_out = {data_in[1087:24],   4'hf,  data_in[23:20],     8'h1,                8'h80};
                    1069: data_out = {data_in[1087:24],   3'h7,  data_in[23:19],     8'h3,                8'h80};
                    1070: data_out = {data_in[1087:24],   2'h3,  data_in[23:18],     8'h7,                8'h80};
                    1071: data_out = {data_in[1087:24],   1'h1,  data_in[23:17],     8'hf,                8'h80};
                    1072: data_out = {data_in[1087:16],                              8'h1f,               8'h80};

                    1073: data_out = {data_in[1087:16],   7'h1f, data_in[15],                             8'h80};
                    1074: data_out = {data_in[1087:16],   6'h1f, data_in[15:14],                          8'h80};
                    1075: data_out = {data_in[1087:16],   5'h1f, data_in[15:13],                          8'h80};
                    1076: data_out = {data_in[1087:16],   4'hf,  data_in[15:12],                          8'h81};
                    1077: data_out = {data_in[1087:16],   3'h7,  data_in[15:11],                          8'h83};
                    1078: data_out = {data_in[1087:16],   2'h3,  data_in[15:10],                          8'h87};
                    1079: data_out = {data_in[1087:16],   1'h1,  data_in[15:9],                           8'h8f};
                    1080: data_out = {data_in[1087:8],                                                    8'h9f};

                    1081: data_out = {data_in[1087:8],    7'h5f, data_in[7]                                    };
                    1082: data_out = {data_in[1087:8],    6'h3f, data_in[7:6]                                  };
						  default: data_out = data_in;
                endcase
                data_next = 1088'b0;
            end
        end else begin
            data_out = data_in;
            data_next = 1088'b0;            
        end
    end

endmodule
